
module mips_16_core_top ( clk, pc );
  output [7:0] pc;
  input clk;
  wire   pipeline_stall_n, branch_taken, reg_write_en, n1, if_stage_inst_n19,
         if_stage_inst_n18, if_stage_inst_n17, if_stage_inst_n16,
         if_stage_inst_n15, if_stage_inst_n14, if_stage_inst_n13,
         if_stage_inst_n12, if_stage_inst_u3_u1_z_7, if_stage_inst_u3_u1_z_4,
         if_stage_inst_u3_u1_z_3, if_stage_inst_u3_u1_z_2,
         if_stage_inst_u3_u1_z_1, if_stage_inst_u3_u1_z_0,
         if_stage_inst_instruction_0_, if_stage_inst_n29, if_stage_inst_n28,
         if_stage_inst_n27, if_stage_inst_n26, if_stage_inst_n25,
         if_stage_inst_n24, if_stage_inst_n23, if_stage_inst_n22,
         if_stage_inst_imem_instruction_15_, if_stage_inst_r301_n1,
         id_stage_inst_n66, id_stage_inst_n46, id_stage_inst_n45,
         id_stage_inst_n44, id_stage_inst_n43, id_stage_inst_n42,
         id_stage_inst_n41, id_stage_inst_n40, id_stage_inst_n39,
         id_stage_inst_n38, id_stage_inst_n37, id_stage_inst_n36,
         id_stage_inst_n35, id_stage_inst_n34, id_stage_inst_n33,
         id_stage_inst_n32, id_stage_inst_n31, id_stage_inst_n30,
         id_stage_inst_n29, id_stage_inst_n28, id_stage_inst_n27,
         id_stage_inst_n26, id_stage_inst_n25, id_stage_inst_n24,
         id_stage_inst_n23, id_stage_inst_n22, id_stage_inst_n21,
         id_stage_inst_n20, id_stage_inst_n19, id_stage_inst_n18,
         id_stage_inst_n17, id_stage_inst_n16, id_stage_inst_n15,
         id_stage_inst_n14, id_stage_inst_n13, id_stage_inst_n12,
         id_stage_inst_n11, id_stage_inst_n10, id_stage_inst_n9,
         id_stage_inst_n8, id_stage_inst_n7, id_stage_inst_n6,
         id_stage_inst_n5, id_stage_inst_n4, id_stage_inst_n3,
         id_stage_inst_n2, id_stage_inst_n1, id_stage_inst_n64,
         id_stage_inst_n63, id_stage_inst_n62, id_stage_inst_n61,
         id_stage_inst_n60, id_stage_inst_n59, id_stage_inst_n58,
         id_stage_inst_n57, id_stage_inst_n56, id_stage_inst_n55,
         id_stage_inst_n54, id_stage_inst_n53, id_stage_inst_n52,
         id_stage_inst_n51, id_stage_inst_n50, id_stage_inst_n49,
         id_stage_inst_write_back_en, id_stage_inst_instruction_reg_9_,
         id_stage_inst_instruction_reg_10_, id_stage_inst_instruction_reg_11_,
         id_stage_inst_instruction_reg_12_, id_stage_inst_instruction_reg_13_,
         id_stage_inst_instruction_reg_14_, id_stage_inst_instruction_reg_15_,
         ex_stage_inst_n40, ex_stage_inst_n39, ex_stage_inst_n38,
         ex_stage_inst_n37, ex_stage_inst_n36, ex_stage_inst_n35,
         ex_stage_inst_n34, ex_stage_inst_n33, ex_stage_inst_n32,
         ex_stage_inst_n31, ex_stage_inst_n30, ex_stage_inst_n29,
         ex_stage_inst_n28, ex_stage_inst_n27, ex_stage_inst_n26,
         ex_stage_inst_n25, ex_stage_inst_n24, ex_stage_inst_n23,
         ex_stage_inst_n22, ex_stage_inst_n21, ex_stage_inst_n20,
         ex_stage_inst_n19, ex_stage_inst_n18, ex_stage_inst_n17,
         ex_stage_inst_n16, ex_stage_inst_n15, ex_stage_inst_n14,
         ex_stage_inst_n13, ex_stage_inst_n12, ex_stage_inst_n11,
         ex_stage_inst_n10, ex_stage_inst_n9, ex_stage_inst_n8,
         ex_stage_inst_n7, ex_stage_inst_n6, ex_stage_inst_n5,
         ex_stage_inst_n4, ex_stage_inst_n3, ex_stage_inst_alu_inst_n209,
         ex_stage_inst_alu_inst_n208, ex_stage_inst_alu_inst_n207,
         ex_stage_inst_alu_inst_n206, ex_stage_inst_alu_inst_n205,
         ex_stage_inst_alu_inst_n204, ex_stage_inst_alu_inst_n203,
         ex_stage_inst_alu_inst_n202, ex_stage_inst_alu_inst_n201,
         ex_stage_inst_alu_inst_n200, ex_stage_inst_alu_inst_n199,
         ex_stage_inst_alu_inst_n198, ex_stage_inst_alu_inst_n197,
         ex_stage_inst_alu_inst_n196, ex_stage_inst_alu_inst_n195,
         ex_stage_inst_alu_inst_n194, ex_stage_inst_alu_inst_n193,
         ex_stage_inst_alu_inst_n192, ex_stage_inst_alu_inst_n191,
         ex_stage_inst_alu_inst_n190, ex_stage_inst_alu_inst_n189,
         ex_stage_inst_alu_inst_n188, ex_stage_inst_alu_inst_n187,
         ex_stage_inst_alu_inst_n186, ex_stage_inst_alu_inst_n185,
         ex_stage_inst_alu_inst_n184, ex_stage_inst_alu_inst_n183,
         ex_stage_inst_alu_inst_n182, ex_stage_inst_alu_inst_n181,
         ex_stage_inst_alu_inst_n180, ex_stage_inst_alu_inst_n179,
         ex_stage_inst_alu_inst_n178, ex_stage_inst_alu_inst_n177,
         ex_stage_inst_alu_inst_n176, ex_stage_inst_alu_inst_n175,
         ex_stage_inst_alu_inst_n174, ex_stage_inst_alu_inst_n173,
         ex_stage_inst_alu_inst_n172, ex_stage_inst_alu_inst_n171,
         ex_stage_inst_alu_inst_n170, ex_stage_inst_alu_inst_n169,
         ex_stage_inst_alu_inst_n168, ex_stage_inst_alu_inst_n167,
         ex_stage_inst_alu_inst_n166, ex_stage_inst_alu_inst_n165,
         ex_stage_inst_alu_inst_n164, ex_stage_inst_alu_inst_n163,
         ex_stage_inst_alu_inst_n162, ex_stage_inst_alu_inst_n161,
         ex_stage_inst_alu_inst_n160, ex_stage_inst_alu_inst_n159,
         ex_stage_inst_alu_inst_n158, ex_stage_inst_alu_inst_n157,
         ex_stage_inst_alu_inst_n156, ex_stage_inst_alu_inst_n155,
         ex_stage_inst_alu_inst_n154, ex_stage_inst_alu_inst_n153,
         ex_stage_inst_alu_inst_n152, ex_stage_inst_alu_inst_n151,
         ex_stage_inst_alu_inst_n150, ex_stage_inst_alu_inst_n149,
         ex_stage_inst_alu_inst_n148, ex_stage_inst_alu_inst_n147,
         ex_stage_inst_alu_inst_n146, ex_stage_inst_alu_inst_n145,
         ex_stage_inst_alu_inst_n144, ex_stage_inst_alu_inst_n143,
         ex_stage_inst_alu_inst_n142, ex_stage_inst_alu_inst_n141,
         ex_stage_inst_alu_inst_n140, ex_stage_inst_alu_inst_n139,
         ex_stage_inst_alu_inst_n138, ex_stage_inst_alu_inst_n137,
         ex_stage_inst_alu_inst_n136, ex_stage_inst_alu_inst_n135,
         ex_stage_inst_alu_inst_n134, ex_stage_inst_alu_inst_n133,
         ex_stage_inst_alu_inst_n132, ex_stage_inst_alu_inst_n131,
         ex_stage_inst_alu_inst_n130, ex_stage_inst_alu_inst_n129,
         ex_stage_inst_alu_inst_n128, ex_stage_inst_alu_inst_n127,
         ex_stage_inst_alu_inst_n126, ex_stage_inst_alu_inst_n125,
         ex_stage_inst_alu_inst_n124, ex_stage_inst_alu_inst_n123,
         ex_stage_inst_alu_inst_n122, ex_stage_inst_alu_inst_n121,
         ex_stage_inst_alu_inst_n120, ex_stage_inst_alu_inst_n119,
         ex_stage_inst_alu_inst_n118, ex_stage_inst_alu_inst_n117,
         ex_stage_inst_alu_inst_n116, ex_stage_inst_alu_inst_n115,
         ex_stage_inst_alu_inst_n114, ex_stage_inst_alu_inst_n113,
         ex_stage_inst_alu_inst_n112, ex_stage_inst_alu_inst_n111,
         ex_stage_inst_alu_inst_n110, ex_stage_inst_alu_inst_n109,
         ex_stage_inst_alu_inst_n108, ex_stage_inst_alu_inst_n107,
         ex_stage_inst_alu_inst_n106, ex_stage_inst_alu_inst_n105,
         ex_stage_inst_alu_inst_n104, ex_stage_inst_alu_inst_n103,
         ex_stage_inst_alu_inst_n102, ex_stage_inst_alu_inst_n101,
         ex_stage_inst_alu_inst_n100, ex_stage_inst_alu_inst_n99,
         ex_stage_inst_alu_inst_n98, ex_stage_inst_alu_inst_n97,
         ex_stage_inst_alu_inst_n96, ex_stage_inst_alu_inst_n95,
         ex_stage_inst_alu_inst_n94, ex_stage_inst_alu_inst_n93,
         ex_stage_inst_alu_inst_n92, ex_stage_inst_alu_inst_n91,
         ex_stage_inst_alu_inst_n90, ex_stage_inst_alu_inst_n89,
         ex_stage_inst_alu_inst_n88, ex_stage_inst_alu_inst_n87,
         ex_stage_inst_alu_inst_n86, ex_stage_inst_alu_inst_n85,
         ex_stage_inst_alu_inst_n84, ex_stage_inst_alu_inst_n83,
         ex_stage_inst_alu_inst_n82, ex_stage_inst_alu_inst_n81,
         ex_stage_inst_alu_inst_n80, ex_stage_inst_alu_inst_n79,
         ex_stage_inst_alu_inst_n78, ex_stage_inst_alu_inst_n77,
         ex_stage_inst_alu_inst_n76, ex_stage_inst_alu_inst_n75,
         ex_stage_inst_alu_inst_n74, ex_stage_inst_alu_inst_n73,
         ex_stage_inst_alu_inst_n72, ex_stage_inst_alu_inst_n71,
         ex_stage_inst_alu_inst_n70, ex_stage_inst_alu_inst_n69,
         ex_stage_inst_alu_inst_n68, ex_stage_inst_alu_inst_n67,
         ex_stage_inst_alu_inst_n66, ex_stage_inst_alu_inst_n65,
         ex_stage_inst_alu_inst_n64, ex_stage_inst_alu_inst_n63,
         ex_stage_inst_alu_inst_n62, ex_stage_inst_alu_inst_n61,
         ex_stage_inst_alu_inst_n60, ex_stage_inst_alu_inst_n59,
         ex_stage_inst_alu_inst_n58, ex_stage_inst_alu_inst_n57,
         ex_stage_inst_alu_inst_n56, ex_stage_inst_alu_inst_n55,
         ex_stage_inst_alu_inst_n54, ex_stage_inst_alu_inst_n53,
         ex_stage_inst_alu_inst_n52, ex_stage_inst_alu_inst_n51,
         ex_stage_inst_alu_inst_n50, ex_stage_inst_alu_inst_n49,
         ex_stage_inst_alu_inst_n48, ex_stage_inst_alu_inst_n47,
         ex_stage_inst_alu_inst_n46, ex_stage_inst_alu_inst_n45,
         ex_stage_inst_alu_inst_n44, ex_stage_inst_alu_inst_n43,
         ex_stage_inst_alu_inst_n42, ex_stage_inst_alu_inst_n41,
         ex_stage_inst_alu_inst_n40, ex_stage_inst_alu_inst_n39,
         ex_stage_inst_alu_inst_n38, ex_stage_inst_alu_inst_n37,
         ex_stage_inst_alu_inst_n36, ex_stage_inst_alu_inst_n35,
         ex_stage_inst_alu_inst_n34, ex_stage_inst_alu_inst_n33,
         ex_stage_inst_alu_inst_n32, ex_stage_inst_alu_inst_n31,
         ex_stage_inst_alu_inst_n30, ex_stage_inst_alu_inst_n29,
         ex_stage_inst_alu_inst_n28, ex_stage_inst_alu_inst_n27,
         ex_stage_inst_alu_inst_n25, ex_stage_inst_alu_inst_n24,
         ex_stage_inst_alu_inst_n23, ex_stage_inst_alu_inst_n22,
         ex_stage_inst_alu_inst_n21, ex_stage_inst_alu_inst_n20,
         ex_stage_inst_alu_inst_n19, ex_stage_inst_alu_inst_n18,
         ex_stage_inst_alu_inst_n17, ex_stage_inst_alu_inst_n16,
         ex_stage_inst_alu_inst_n15, ex_stage_inst_alu_inst_n14,
         ex_stage_inst_alu_inst_n13, ex_stage_inst_alu_inst_n12,
         ex_stage_inst_alu_inst_n11, ex_stage_inst_alu_inst_n10,
         ex_stage_inst_alu_inst_n9, ex_stage_inst_alu_inst_n8,
         ex_stage_inst_alu_inst_n7, ex_stage_inst_alu_inst_n6,
         ex_stage_inst_alu_inst_n5, ex_stage_inst_alu_inst_n4,
         ex_stage_inst_alu_inst_n3, ex_stage_inst_alu_inst_n2,
         ex_stage_inst_alu_inst_n1, ex_stage_inst_alu_inst_n26,
         ex_stage_inst_alu_inst_n1600, ex_stage_inst_alu_inst_n1590,
         ex_stage_inst_alu_inst_n1580, ex_stage_inst_alu_inst_n1570,
         ex_stage_inst_alu_inst_n1560, ex_stage_inst_alu_inst_n1550,
         ex_stage_inst_alu_inst_n1540, ex_stage_inst_alu_inst_n1530,
         ex_stage_inst_alu_inst_n1520, ex_stage_inst_alu_inst_n1510,
         ex_stage_inst_alu_inst_n1500, ex_stage_inst_alu_inst_n1490,
         ex_stage_inst_alu_inst_n1480, ex_stage_inst_alu_inst_n1470,
         ex_stage_inst_alu_inst_n1460, ex_stage_inst_alu_inst_n1450,
         ex_stage_inst_alu_inst_n1280, ex_stage_inst_alu_inst_n1270,
         ex_stage_inst_alu_inst_n1260, ex_stage_inst_alu_inst_n1250,
         ex_stage_inst_alu_inst_n1240, ex_stage_inst_alu_inst_n1230,
         ex_stage_inst_alu_inst_n1220, ex_stage_inst_alu_inst_n1210,
         ex_stage_inst_alu_inst_n1200, ex_stage_inst_alu_inst_n1190,
         ex_stage_inst_alu_inst_n1180, ex_stage_inst_alu_inst_n1170,
         ex_stage_inst_alu_inst_n1160, ex_stage_inst_alu_inst_n1150,
         ex_stage_inst_alu_inst_n1140, ex_stage_inst_alu_inst_n1130,
         ex_stage_inst_alu_inst_n640, ex_stage_inst_alu_inst_n630,
         ex_stage_inst_alu_inst_n620, ex_stage_inst_alu_inst_n610,
         ex_stage_inst_alu_inst_n600, ex_stage_inst_alu_inst_n590,
         ex_stage_inst_alu_inst_n580, ex_stage_inst_alu_inst_n570,
         ex_stage_inst_alu_inst_n560, ex_stage_inst_alu_inst_n550,
         ex_stage_inst_alu_inst_n540, ex_stage_inst_alu_inst_n530,
         ex_stage_inst_alu_inst_n520, ex_stage_inst_alu_inst_n510,
         ex_stage_inst_alu_inst_n500, ex_stage_inst_alu_inst_n490,
         ex_stage_inst_alu_inst_r316_carry_1_,
         ex_stage_inst_alu_inst_r316_carry_2_,
         ex_stage_inst_alu_inst_r316_carry_3_,
         ex_stage_inst_alu_inst_r316_carry_4_,
         ex_stage_inst_alu_inst_r316_carry_5_,
         ex_stage_inst_alu_inst_r316_carry_6_,
         ex_stage_inst_alu_inst_r316_carry_7_,
         ex_stage_inst_alu_inst_r316_carry_8_,
         ex_stage_inst_alu_inst_r316_carry_9_,
         ex_stage_inst_alu_inst_r316_carry_10_,
         ex_stage_inst_alu_inst_r316_carry_11_,
         ex_stage_inst_alu_inst_r316_carry_12_,
         ex_stage_inst_alu_inst_r316_carry_13_,
         ex_stage_inst_alu_inst_r316_carry_14_,
         ex_stage_inst_alu_inst_r316_carry_15_,
         ex_stage_inst_alu_inst_sll_36_n146,
         ex_stage_inst_alu_inst_sll_36_n145, ex_stage_inst_alu_inst_sll_36_n91,
         ex_stage_inst_alu_inst_sll_36_n89, ex_stage_inst_alu_inst_sll_36_n88,
         ex_stage_inst_alu_inst_sll_36_n87, ex_stage_inst_alu_inst_sll_36_n86,
         ex_stage_inst_alu_inst_sll_36_n85, ex_stage_inst_alu_inst_sll_36_n84,
         ex_stage_inst_alu_inst_sll_36_n82, ex_stage_inst_alu_inst_sll_36_n81,
         ex_stage_inst_alu_inst_sll_36_n80, ex_stage_inst_alu_inst_sll_36_n79,
         ex_stage_inst_alu_inst_sll_36_n78, ex_stage_inst_alu_inst_sll_36_n77,
         ex_stage_inst_alu_inst_sll_36_n76, ex_stage_inst_alu_inst_sll_36_n75,
         ex_stage_inst_alu_inst_sll_36_n74, ex_stage_inst_alu_inst_sll_36_n73,
         ex_stage_inst_alu_inst_sll_36_n72, ex_stage_inst_alu_inst_sll_36_n71,
         ex_stage_inst_alu_inst_sll_36_n70, ex_stage_inst_alu_inst_sll_36_n69,
         ex_stage_inst_alu_inst_sll_36_n68, ex_stage_inst_alu_inst_sll_36_n67,
         ex_stage_inst_alu_inst_sll_36_n66, ex_stage_inst_alu_inst_sll_36_n65,
         ex_stage_inst_alu_inst_sll_36_n64, ex_stage_inst_alu_inst_sll_36_n63,
         ex_stage_inst_alu_inst_sll_36_n62, ex_stage_inst_alu_inst_sll_36_n61,
         ex_stage_inst_alu_inst_sll_36_n60, ex_stage_inst_alu_inst_sll_36_n59,
         ex_stage_inst_alu_inst_sll_36_n58, ex_stage_inst_alu_inst_sll_36_n57,
         ex_stage_inst_alu_inst_sll_36_n56, ex_stage_inst_alu_inst_sll_36_n55,
         ex_stage_inst_alu_inst_sll_36_n54, ex_stage_inst_alu_inst_sll_36_n53,
         ex_stage_inst_alu_inst_sll_36_n52, ex_stage_inst_alu_inst_sll_36_n51,
         ex_stage_inst_alu_inst_sll_36_n50, ex_stage_inst_alu_inst_sll_36_n49,
         ex_stage_inst_alu_inst_sll_36_n48, ex_stage_inst_alu_inst_sll_36_n47,
         ex_stage_inst_alu_inst_sll_36_n46, ex_stage_inst_alu_inst_sll_36_n45,
         ex_stage_inst_alu_inst_sll_36_n44, ex_stage_inst_alu_inst_sll_36_n43,
         ex_stage_inst_alu_inst_sll_36_n42, ex_stage_inst_alu_inst_sll_36_n41,
         ex_stage_inst_alu_inst_sll_36_n40, ex_stage_inst_alu_inst_sll_36_n39,
         ex_stage_inst_alu_inst_sll_36_n38, ex_stage_inst_alu_inst_sll_36_n37,
         ex_stage_inst_alu_inst_sll_36_n36, ex_stage_inst_alu_inst_sll_36_n35,
         ex_stage_inst_alu_inst_sll_36_n34, ex_stage_inst_alu_inst_sll_36_n33,
         ex_stage_inst_alu_inst_sll_36_n32, ex_stage_inst_alu_inst_sll_36_n31,
         ex_stage_inst_alu_inst_sll_36_n30, ex_stage_inst_alu_inst_sll_36_n29,
         ex_stage_inst_alu_inst_sll_36_n28, ex_stage_inst_alu_inst_sll_36_n27,
         ex_stage_inst_alu_inst_sll_36_n26, ex_stage_inst_alu_inst_sll_36_n25,
         ex_stage_inst_alu_inst_sll_36_n24, ex_stage_inst_alu_inst_sll_36_n23,
         ex_stage_inst_alu_inst_sll_36_n22, ex_stage_inst_alu_inst_sll_36_n21,
         ex_stage_inst_alu_inst_sll_36_n20, ex_stage_inst_alu_inst_sll_36_n19,
         ex_stage_inst_alu_inst_sll_36_n18, ex_stage_inst_alu_inst_sll_36_n17,
         ex_stage_inst_alu_inst_sll_36_n16, ex_stage_inst_alu_inst_sll_36_n15,
         ex_stage_inst_alu_inst_sll_36_n14, ex_stage_inst_alu_inst_sll_36_n13,
         ex_stage_inst_alu_inst_sll_36_n12, ex_stage_inst_alu_inst_sll_36_n11,
         ex_stage_inst_alu_inst_sll_36_n10, ex_stage_inst_alu_inst_sll_36_n9,
         ex_stage_inst_alu_inst_sll_36_n8, ex_stage_inst_alu_inst_sll_36_n7,
         ex_stage_inst_alu_inst_sll_36_n6, ex_stage_inst_alu_inst_sll_36_n5,
         ex_stage_inst_alu_inst_sll_36_n4, ex_stage_inst_alu_inst_sll_36_n3,
         ex_stage_inst_alu_inst_sll_36_n2, ex_stage_inst_alu_inst_srl_40_n148,
         ex_stage_inst_alu_inst_srl_40_n147, ex_stage_inst_alu_inst_srl_40_n91,
         ex_stage_inst_alu_inst_srl_40_n89, ex_stage_inst_alu_inst_srl_40_n88,
         ex_stage_inst_alu_inst_srl_40_n87, ex_stage_inst_alu_inst_srl_40_n86,
         ex_stage_inst_alu_inst_srl_40_n85, ex_stage_inst_alu_inst_srl_40_n84,
         ex_stage_inst_alu_inst_srl_40_n82, ex_stage_inst_alu_inst_srl_40_n81,
         ex_stage_inst_alu_inst_srl_40_n80, ex_stage_inst_alu_inst_srl_40_n79,
         ex_stage_inst_alu_inst_srl_40_n78, ex_stage_inst_alu_inst_srl_40_n77,
         ex_stage_inst_alu_inst_srl_40_n76, ex_stage_inst_alu_inst_srl_40_n75,
         ex_stage_inst_alu_inst_srl_40_n74, ex_stage_inst_alu_inst_srl_40_n73,
         ex_stage_inst_alu_inst_srl_40_n72, ex_stage_inst_alu_inst_srl_40_n71,
         ex_stage_inst_alu_inst_srl_40_n70, ex_stage_inst_alu_inst_srl_40_n69,
         ex_stage_inst_alu_inst_srl_40_n68, ex_stage_inst_alu_inst_srl_40_n67,
         ex_stage_inst_alu_inst_srl_40_n66, ex_stage_inst_alu_inst_srl_40_n65,
         ex_stage_inst_alu_inst_srl_40_n64, ex_stage_inst_alu_inst_srl_40_n63,
         ex_stage_inst_alu_inst_srl_40_n62, ex_stage_inst_alu_inst_srl_40_n61,
         ex_stage_inst_alu_inst_srl_40_n60, ex_stage_inst_alu_inst_srl_40_n59,
         ex_stage_inst_alu_inst_srl_40_n58, ex_stage_inst_alu_inst_srl_40_n57,
         ex_stage_inst_alu_inst_srl_40_n56, ex_stage_inst_alu_inst_srl_40_n55,
         ex_stage_inst_alu_inst_srl_40_n54, ex_stage_inst_alu_inst_srl_40_n53,
         ex_stage_inst_alu_inst_srl_40_n52, ex_stage_inst_alu_inst_srl_40_n51,
         ex_stage_inst_alu_inst_srl_40_n50, ex_stage_inst_alu_inst_srl_40_n49,
         ex_stage_inst_alu_inst_srl_40_n48, ex_stage_inst_alu_inst_srl_40_n47,
         ex_stage_inst_alu_inst_srl_40_n46, ex_stage_inst_alu_inst_srl_40_n45,
         ex_stage_inst_alu_inst_srl_40_n44, ex_stage_inst_alu_inst_srl_40_n43,
         ex_stage_inst_alu_inst_srl_40_n42, ex_stage_inst_alu_inst_srl_40_n41,
         ex_stage_inst_alu_inst_srl_40_n40, ex_stage_inst_alu_inst_srl_40_n39,
         ex_stage_inst_alu_inst_srl_40_n38, ex_stage_inst_alu_inst_srl_40_n37,
         ex_stage_inst_alu_inst_srl_40_n36, ex_stage_inst_alu_inst_srl_40_n35,
         ex_stage_inst_alu_inst_srl_40_n34, ex_stage_inst_alu_inst_srl_40_n33,
         ex_stage_inst_alu_inst_srl_40_n32, ex_stage_inst_alu_inst_srl_40_n31,
         ex_stage_inst_alu_inst_srl_40_n30, ex_stage_inst_alu_inst_srl_40_n29,
         ex_stage_inst_alu_inst_srl_40_n28, ex_stage_inst_alu_inst_srl_40_n27,
         ex_stage_inst_alu_inst_srl_40_n26, ex_stage_inst_alu_inst_srl_40_n25,
         ex_stage_inst_alu_inst_srl_40_n24, ex_stage_inst_alu_inst_srl_40_n23,
         ex_stage_inst_alu_inst_srl_40_n22, ex_stage_inst_alu_inst_srl_40_n21,
         ex_stage_inst_alu_inst_srl_40_n20, ex_stage_inst_alu_inst_srl_40_n19,
         ex_stage_inst_alu_inst_srl_40_n18, ex_stage_inst_alu_inst_srl_40_n17,
         ex_stage_inst_alu_inst_srl_40_n16, ex_stage_inst_alu_inst_srl_40_n15,
         ex_stage_inst_alu_inst_srl_40_n14, ex_stage_inst_alu_inst_srl_40_n13,
         ex_stage_inst_alu_inst_srl_40_n12, ex_stage_inst_alu_inst_srl_40_n11,
         ex_stage_inst_alu_inst_srl_40_n10, ex_stage_inst_alu_inst_srl_40_n9,
         ex_stage_inst_alu_inst_srl_40_n8, ex_stage_inst_alu_inst_srl_40_n7,
         ex_stage_inst_alu_inst_srl_40_n6, ex_stage_inst_alu_inst_srl_40_n5,
         ex_stage_inst_alu_inst_srl_40_n4, ex_stage_inst_alu_inst_srl_40_n3,
         ex_stage_inst_alu_inst_srl_40_n2, mem_stage_inst_n39,
         mem_stage_inst_n38, mem_stage_inst_n37, mem_stage_inst_n36,
         mem_stage_inst_n35, mem_stage_inst_n34, mem_stage_inst_n33,
         mem_stage_inst_n32, mem_stage_inst_n31, mem_stage_inst_n30,
         mem_stage_inst_n29, mem_stage_inst_n28, mem_stage_inst_n27,
         mem_stage_inst_n26, mem_stage_inst_n25, mem_stage_inst_n24,
         mem_stage_inst_n23, mem_stage_inst_n22, mem_stage_inst_n21,
         mem_stage_inst_n20, mem_stage_inst_n19, mem_stage_inst_n18,
         mem_stage_inst_n17, mem_stage_inst_n16, mem_stage_inst_n15,
         mem_stage_inst_n14, mem_stage_inst_n13, mem_stage_inst_n12,
         mem_stage_inst_n11, mem_stage_inst_n10, mem_stage_inst_n9,
         mem_stage_inst_n8, mem_stage_inst_n7, mem_stage_inst_n6,
         mem_stage_inst_n5, mem_stage_inst_n4, mem_stage_inst_n3,
         mem_stage_inst_dmem_n5969, mem_stage_inst_dmem_n5968,
         mem_stage_inst_dmem_n5967, mem_stage_inst_dmem_n5966,
         mem_stage_inst_dmem_n5965, mem_stage_inst_dmem_n5964,
         mem_stage_inst_dmem_n5963, mem_stage_inst_dmem_n5962,
         mem_stage_inst_dmem_n5961, mem_stage_inst_dmem_n5960,
         mem_stage_inst_dmem_n5959, mem_stage_inst_dmem_n5958,
         mem_stage_inst_dmem_n5957, mem_stage_inst_dmem_n5956,
         mem_stage_inst_dmem_n5955, mem_stage_inst_dmem_n5954,
         mem_stage_inst_dmem_n5953, mem_stage_inst_dmem_n5952,
         mem_stage_inst_dmem_n5951, mem_stage_inst_dmem_n5950,
         mem_stage_inst_dmem_n5949, mem_stage_inst_dmem_n5948,
         mem_stage_inst_dmem_n5947, mem_stage_inst_dmem_n5946,
         mem_stage_inst_dmem_n5945, mem_stage_inst_dmem_n5944,
         mem_stage_inst_dmem_n5943, mem_stage_inst_dmem_n5942,
         mem_stage_inst_dmem_n5941, mem_stage_inst_dmem_n5940,
         mem_stage_inst_dmem_n5939, mem_stage_inst_dmem_n5938,
         mem_stage_inst_dmem_n5937, mem_stage_inst_dmem_n5936,
         mem_stage_inst_dmem_n5935, mem_stage_inst_dmem_n5934,
         mem_stage_inst_dmem_n5933, mem_stage_inst_dmem_n5932,
         mem_stage_inst_dmem_n5931, mem_stage_inst_dmem_n5930,
         mem_stage_inst_dmem_n5929, mem_stage_inst_dmem_n5928,
         mem_stage_inst_dmem_n5927, mem_stage_inst_dmem_n5926,
         mem_stage_inst_dmem_n5925, mem_stage_inst_dmem_n5924,
         mem_stage_inst_dmem_n5923, mem_stage_inst_dmem_n5922,
         mem_stage_inst_dmem_n5921, mem_stage_inst_dmem_n5920,
         mem_stage_inst_dmem_n5919, mem_stage_inst_dmem_n5918,
         mem_stage_inst_dmem_n5917, mem_stage_inst_dmem_n5916,
         mem_stage_inst_dmem_n5915, mem_stage_inst_dmem_n5914,
         mem_stage_inst_dmem_n5913, mem_stage_inst_dmem_n5912,
         mem_stage_inst_dmem_n5911, mem_stage_inst_dmem_n5910,
         mem_stage_inst_dmem_n5909, mem_stage_inst_dmem_n5908,
         mem_stage_inst_dmem_n5907, mem_stage_inst_dmem_n5906,
         mem_stage_inst_dmem_n5905, mem_stage_inst_dmem_n5904,
         mem_stage_inst_dmem_n5903, mem_stage_inst_dmem_n5902,
         mem_stage_inst_dmem_n5901, mem_stage_inst_dmem_n5900,
         mem_stage_inst_dmem_n5899, mem_stage_inst_dmem_n5898,
         mem_stage_inst_dmem_n5897, mem_stage_inst_dmem_n5896,
         mem_stage_inst_dmem_n5895, mem_stage_inst_dmem_n5894,
         mem_stage_inst_dmem_n5893, mem_stage_inst_dmem_n5892,
         mem_stage_inst_dmem_n5891, mem_stage_inst_dmem_n5890,
         mem_stage_inst_dmem_n5889, mem_stage_inst_dmem_n5888,
         mem_stage_inst_dmem_n5887, mem_stage_inst_dmem_n5886,
         mem_stage_inst_dmem_n5885, mem_stage_inst_dmem_n5884,
         mem_stage_inst_dmem_n5883, mem_stage_inst_dmem_n5882,
         mem_stage_inst_dmem_n5881, mem_stage_inst_dmem_n5880,
         mem_stage_inst_dmem_n5879, mem_stage_inst_dmem_n5878,
         mem_stage_inst_dmem_n5877, mem_stage_inst_dmem_n5876,
         mem_stage_inst_dmem_n5875, mem_stage_inst_dmem_n5874,
         mem_stage_inst_dmem_n5873, mem_stage_inst_dmem_n5872,
         mem_stage_inst_dmem_n5871, mem_stage_inst_dmem_n5870,
         mem_stage_inst_dmem_n5869, mem_stage_inst_dmem_n5868,
         mem_stage_inst_dmem_n5867, mem_stage_inst_dmem_n5866,
         mem_stage_inst_dmem_n5865, mem_stage_inst_dmem_n5864,
         mem_stage_inst_dmem_n5863, mem_stage_inst_dmem_n5862,
         mem_stage_inst_dmem_n5861, mem_stage_inst_dmem_n5860,
         mem_stage_inst_dmem_n5859, mem_stage_inst_dmem_n5858,
         mem_stage_inst_dmem_n5857, mem_stage_inst_dmem_n5856,
         mem_stage_inst_dmem_n5855, mem_stage_inst_dmem_n5854,
         mem_stage_inst_dmem_n5853, mem_stage_inst_dmem_n5852,
         mem_stage_inst_dmem_n5851, mem_stage_inst_dmem_n5850,
         mem_stage_inst_dmem_n5849, mem_stage_inst_dmem_n5848,
         mem_stage_inst_dmem_n5847, mem_stage_inst_dmem_n5846,
         mem_stage_inst_dmem_n5845, mem_stage_inst_dmem_n5844,
         mem_stage_inst_dmem_n5843, mem_stage_inst_dmem_n5842,
         mem_stage_inst_dmem_n5841, mem_stage_inst_dmem_n5840,
         mem_stage_inst_dmem_n5839, mem_stage_inst_dmem_n5838,
         mem_stage_inst_dmem_n5837, mem_stage_inst_dmem_n5836,
         mem_stage_inst_dmem_n5835, mem_stage_inst_dmem_n5834,
         mem_stage_inst_dmem_n5833, mem_stage_inst_dmem_n5832,
         mem_stage_inst_dmem_n5831, mem_stage_inst_dmem_n5830,
         mem_stage_inst_dmem_n5829, mem_stage_inst_dmem_n5828,
         mem_stage_inst_dmem_n5827, mem_stage_inst_dmem_n5826,
         mem_stage_inst_dmem_n5825, mem_stage_inst_dmem_n5824,
         mem_stage_inst_dmem_n5823, mem_stage_inst_dmem_n5822,
         mem_stage_inst_dmem_n5821, mem_stage_inst_dmem_n5820,
         mem_stage_inst_dmem_n5819, mem_stage_inst_dmem_n5818,
         mem_stage_inst_dmem_n5817, mem_stage_inst_dmem_n5816,
         mem_stage_inst_dmem_n5815, mem_stage_inst_dmem_n5814,
         mem_stage_inst_dmem_n5813, mem_stage_inst_dmem_n5812,
         mem_stage_inst_dmem_n5811, mem_stage_inst_dmem_n5810,
         mem_stage_inst_dmem_n5809, mem_stage_inst_dmem_n5808,
         mem_stage_inst_dmem_n5807, mem_stage_inst_dmem_n5806,
         mem_stage_inst_dmem_n5805, mem_stage_inst_dmem_n5804,
         mem_stage_inst_dmem_n5803, mem_stage_inst_dmem_n5802,
         mem_stage_inst_dmem_n5801, mem_stage_inst_dmem_n5800,
         mem_stage_inst_dmem_n5799, mem_stage_inst_dmem_n5798,
         mem_stage_inst_dmem_n5797, mem_stage_inst_dmem_n5796,
         mem_stage_inst_dmem_n5795, mem_stage_inst_dmem_n5794,
         mem_stage_inst_dmem_n5793, mem_stage_inst_dmem_n5792,
         mem_stage_inst_dmem_n5791, mem_stage_inst_dmem_n5790,
         mem_stage_inst_dmem_n5789, mem_stage_inst_dmem_n5788,
         mem_stage_inst_dmem_n5787, mem_stage_inst_dmem_n5786,
         mem_stage_inst_dmem_n5785, mem_stage_inst_dmem_n5784,
         mem_stage_inst_dmem_n5783, mem_stage_inst_dmem_n5782,
         mem_stage_inst_dmem_n5781, mem_stage_inst_dmem_n5780,
         mem_stage_inst_dmem_n5779, mem_stage_inst_dmem_n5778,
         mem_stage_inst_dmem_n5777, mem_stage_inst_dmem_n5776,
         mem_stage_inst_dmem_n5775, mem_stage_inst_dmem_n5774,
         mem_stage_inst_dmem_n5773, mem_stage_inst_dmem_n5772,
         mem_stage_inst_dmem_n5771, mem_stage_inst_dmem_n5770,
         mem_stage_inst_dmem_n5769, mem_stage_inst_dmem_n5768,
         mem_stage_inst_dmem_n5767, mem_stage_inst_dmem_n5766,
         mem_stage_inst_dmem_n5765, mem_stage_inst_dmem_n5764,
         mem_stage_inst_dmem_n5763, mem_stage_inst_dmem_n5762,
         mem_stage_inst_dmem_n5761, mem_stage_inst_dmem_n5760,
         mem_stage_inst_dmem_n5759, mem_stage_inst_dmem_n5758,
         mem_stage_inst_dmem_n5757, mem_stage_inst_dmem_n5756,
         mem_stage_inst_dmem_n5755, mem_stage_inst_dmem_n5754,
         mem_stage_inst_dmem_n5753, mem_stage_inst_dmem_n5752,
         mem_stage_inst_dmem_n5751, mem_stage_inst_dmem_n5750,
         mem_stage_inst_dmem_n5749, mem_stage_inst_dmem_n5748,
         mem_stage_inst_dmem_n5747, mem_stage_inst_dmem_n5746,
         mem_stage_inst_dmem_n5745, mem_stage_inst_dmem_n5744,
         mem_stage_inst_dmem_n5743, mem_stage_inst_dmem_n5742,
         mem_stage_inst_dmem_n5741, mem_stage_inst_dmem_n5740,
         mem_stage_inst_dmem_n5739, mem_stage_inst_dmem_n5738,
         mem_stage_inst_dmem_n5737, mem_stage_inst_dmem_n5736,
         mem_stage_inst_dmem_n5735, mem_stage_inst_dmem_n5734,
         mem_stage_inst_dmem_n5733, mem_stage_inst_dmem_n5732,
         mem_stage_inst_dmem_n5731, mem_stage_inst_dmem_n5730,
         mem_stage_inst_dmem_n5729, mem_stage_inst_dmem_n5728,
         mem_stage_inst_dmem_n5727, mem_stage_inst_dmem_n5726,
         mem_stage_inst_dmem_n5725, mem_stage_inst_dmem_n5724,
         mem_stage_inst_dmem_n5723, mem_stage_inst_dmem_n5722,
         mem_stage_inst_dmem_n5721, mem_stage_inst_dmem_n5720,
         mem_stage_inst_dmem_n5719, mem_stage_inst_dmem_n5718,
         mem_stage_inst_dmem_n5717, mem_stage_inst_dmem_n5716,
         mem_stage_inst_dmem_n5715, mem_stage_inst_dmem_n5714,
         mem_stage_inst_dmem_n5713, mem_stage_inst_dmem_n5712,
         mem_stage_inst_dmem_n5711, mem_stage_inst_dmem_n5710,
         mem_stage_inst_dmem_n5709, mem_stage_inst_dmem_n5708,
         mem_stage_inst_dmem_n5707, mem_stage_inst_dmem_n5706,
         mem_stage_inst_dmem_n5705, mem_stage_inst_dmem_n5704,
         mem_stage_inst_dmem_n5703, mem_stage_inst_dmem_n5702,
         mem_stage_inst_dmem_n5701, mem_stage_inst_dmem_n5700,
         mem_stage_inst_dmem_n5699, mem_stage_inst_dmem_n5698,
         mem_stage_inst_dmem_n5697, mem_stage_inst_dmem_n5696,
         mem_stage_inst_dmem_n5695, mem_stage_inst_dmem_n5694,
         mem_stage_inst_dmem_n5693, mem_stage_inst_dmem_n5692,
         mem_stage_inst_dmem_n5691, mem_stage_inst_dmem_n5690,
         mem_stage_inst_dmem_n5689, mem_stage_inst_dmem_n5688,
         mem_stage_inst_dmem_n5687, mem_stage_inst_dmem_n5686,
         mem_stage_inst_dmem_n5685, mem_stage_inst_dmem_n5684,
         mem_stage_inst_dmem_n5683, mem_stage_inst_dmem_n5682,
         mem_stage_inst_dmem_n5681, mem_stage_inst_dmem_n5680,
         mem_stage_inst_dmem_n5679, mem_stage_inst_dmem_n5678,
         mem_stage_inst_dmem_n5677, mem_stage_inst_dmem_n5676,
         mem_stage_inst_dmem_n5675, mem_stage_inst_dmem_n5674,
         mem_stage_inst_dmem_n5673, mem_stage_inst_dmem_n5672,
         mem_stage_inst_dmem_n5671, mem_stage_inst_dmem_n5670,
         mem_stage_inst_dmem_n5669, mem_stage_inst_dmem_n5668,
         mem_stage_inst_dmem_n5667, mem_stage_inst_dmem_n5666,
         mem_stage_inst_dmem_n5665, mem_stage_inst_dmem_n5664,
         mem_stage_inst_dmem_n5663, mem_stage_inst_dmem_n5662,
         mem_stage_inst_dmem_n5661, mem_stage_inst_dmem_n5660,
         mem_stage_inst_dmem_n5659, mem_stage_inst_dmem_n5658,
         mem_stage_inst_dmem_n5657, mem_stage_inst_dmem_n5656,
         mem_stage_inst_dmem_n5655, mem_stage_inst_dmem_n5654,
         mem_stage_inst_dmem_n5653, mem_stage_inst_dmem_n5652,
         mem_stage_inst_dmem_n5651, mem_stage_inst_dmem_n5650,
         mem_stage_inst_dmem_n5649, mem_stage_inst_dmem_n5648,
         mem_stage_inst_dmem_n5647, mem_stage_inst_dmem_n5646,
         mem_stage_inst_dmem_n5645, mem_stage_inst_dmem_n5644,
         mem_stage_inst_dmem_n5643, mem_stage_inst_dmem_n5642,
         mem_stage_inst_dmem_n5641, mem_stage_inst_dmem_n5640,
         mem_stage_inst_dmem_n5639, mem_stage_inst_dmem_n5638,
         mem_stage_inst_dmem_n5637, mem_stage_inst_dmem_n5636,
         mem_stage_inst_dmem_n5635, mem_stage_inst_dmem_n5634,
         mem_stage_inst_dmem_n5633, mem_stage_inst_dmem_n5632,
         mem_stage_inst_dmem_n5631, mem_stage_inst_dmem_n5630,
         mem_stage_inst_dmem_n5629, mem_stage_inst_dmem_n5628,
         mem_stage_inst_dmem_n5627, mem_stage_inst_dmem_n5626,
         mem_stage_inst_dmem_n5625, mem_stage_inst_dmem_n5624,
         mem_stage_inst_dmem_n5623, mem_stage_inst_dmem_n5622,
         mem_stage_inst_dmem_n5621, mem_stage_inst_dmem_n5620,
         mem_stage_inst_dmem_n5619, mem_stage_inst_dmem_n5618,
         mem_stage_inst_dmem_n5617, mem_stage_inst_dmem_n5616,
         mem_stage_inst_dmem_n5615, mem_stage_inst_dmem_n5614,
         mem_stage_inst_dmem_n5613, mem_stage_inst_dmem_n5612,
         mem_stage_inst_dmem_n5611, mem_stage_inst_dmem_n5610,
         mem_stage_inst_dmem_n5609, mem_stage_inst_dmem_n5608,
         mem_stage_inst_dmem_n5607, mem_stage_inst_dmem_n5606,
         mem_stage_inst_dmem_n5605, mem_stage_inst_dmem_n5604,
         mem_stage_inst_dmem_n5603, mem_stage_inst_dmem_n5602,
         mem_stage_inst_dmem_n5601, mem_stage_inst_dmem_n5600,
         mem_stage_inst_dmem_n5599, mem_stage_inst_dmem_n5598,
         mem_stage_inst_dmem_n5597, mem_stage_inst_dmem_n5596,
         mem_stage_inst_dmem_n5595, mem_stage_inst_dmem_n5594,
         mem_stage_inst_dmem_n5593, mem_stage_inst_dmem_n5592,
         mem_stage_inst_dmem_n5591, mem_stage_inst_dmem_n5590,
         mem_stage_inst_dmem_n5589, mem_stage_inst_dmem_n5588,
         mem_stage_inst_dmem_n5587, mem_stage_inst_dmem_n5586,
         mem_stage_inst_dmem_n5585, mem_stage_inst_dmem_n5584,
         mem_stage_inst_dmem_n5583, mem_stage_inst_dmem_n5582,
         mem_stage_inst_dmem_n5581, mem_stage_inst_dmem_n5580,
         mem_stage_inst_dmem_n5579, mem_stage_inst_dmem_n5578,
         mem_stage_inst_dmem_n5577, mem_stage_inst_dmem_n5576,
         mem_stage_inst_dmem_n5575, mem_stage_inst_dmem_n5574,
         mem_stage_inst_dmem_n5573, mem_stage_inst_dmem_n5572,
         mem_stage_inst_dmem_n5571, mem_stage_inst_dmem_n5570,
         mem_stage_inst_dmem_n5569, mem_stage_inst_dmem_n5568,
         mem_stage_inst_dmem_n5567, mem_stage_inst_dmem_n5566,
         mem_stage_inst_dmem_n5565, mem_stage_inst_dmem_n5564,
         mem_stage_inst_dmem_n5563, mem_stage_inst_dmem_n5562,
         mem_stage_inst_dmem_n5561, mem_stage_inst_dmem_n5560,
         mem_stage_inst_dmem_n5559, mem_stage_inst_dmem_n5558,
         mem_stage_inst_dmem_n5557, mem_stage_inst_dmem_n5556,
         mem_stage_inst_dmem_n5555, mem_stage_inst_dmem_n5554,
         mem_stage_inst_dmem_n5553, mem_stage_inst_dmem_n5552,
         mem_stage_inst_dmem_n5551, mem_stage_inst_dmem_n5550,
         mem_stage_inst_dmem_n5549, mem_stage_inst_dmem_n5548,
         mem_stage_inst_dmem_n5547, mem_stage_inst_dmem_n5546,
         mem_stage_inst_dmem_n5545, mem_stage_inst_dmem_n5544,
         mem_stage_inst_dmem_n5543, mem_stage_inst_dmem_n5542,
         mem_stage_inst_dmem_n5541, mem_stage_inst_dmem_n5540,
         mem_stage_inst_dmem_n5539, mem_stage_inst_dmem_n5538,
         mem_stage_inst_dmem_n5537, mem_stage_inst_dmem_n5536,
         mem_stage_inst_dmem_n5535, mem_stage_inst_dmem_n5534,
         mem_stage_inst_dmem_n5533, mem_stage_inst_dmem_n5532,
         mem_stage_inst_dmem_n5531, mem_stage_inst_dmem_n5530,
         mem_stage_inst_dmem_n5529, mem_stage_inst_dmem_n5528,
         mem_stage_inst_dmem_n5527, mem_stage_inst_dmem_n5526,
         mem_stage_inst_dmem_n5525, mem_stage_inst_dmem_n5524,
         mem_stage_inst_dmem_n5523, mem_stage_inst_dmem_n5522,
         mem_stage_inst_dmem_n5521, mem_stage_inst_dmem_n5520,
         mem_stage_inst_dmem_n5519, mem_stage_inst_dmem_n5518,
         mem_stage_inst_dmem_n5517, mem_stage_inst_dmem_n5516,
         mem_stage_inst_dmem_n5515, mem_stage_inst_dmem_n5514,
         mem_stage_inst_dmem_n5513, mem_stage_inst_dmem_n5512,
         mem_stage_inst_dmem_n5511, mem_stage_inst_dmem_n5510,
         mem_stage_inst_dmem_n5509, mem_stage_inst_dmem_n5508,
         mem_stage_inst_dmem_n5507, mem_stage_inst_dmem_n5506,
         mem_stage_inst_dmem_n5505, mem_stage_inst_dmem_n5504,
         mem_stage_inst_dmem_n5503, mem_stage_inst_dmem_n5502,
         mem_stage_inst_dmem_n5501, mem_stage_inst_dmem_n5500,
         mem_stage_inst_dmem_n5499, mem_stage_inst_dmem_n5498,
         mem_stage_inst_dmem_n5497, mem_stage_inst_dmem_n5496,
         mem_stage_inst_dmem_n5495, mem_stage_inst_dmem_n5494,
         mem_stage_inst_dmem_n5493, mem_stage_inst_dmem_n5492,
         mem_stage_inst_dmem_n5491, mem_stage_inst_dmem_n5490,
         mem_stage_inst_dmem_n5489, mem_stage_inst_dmem_n5488,
         mem_stage_inst_dmem_n5487, mem_stage_inst_dmem_n5486,
         mem_stage_inst_dmem_n5485, mem_stage_inst_dmem_n5484,
         mem_stage_inst_dmem_n5483, mem_stage_inst_dmem_n5482,
         mem_stage_inst_dmem_n5481, mem_stage_inst_dmem_n5480,
         mem_stage_inst_dmem_n5479, mem_stage_inst_dmem_n5478,
         mem_stage_inst_dmem_n5477, mem_stage_inst_dmem_n5476,
         mem_stage_inst_dmem_n5475, mem_stage_inst_dmem_n5474,
         mem_stage_inst_dmem_n5473, mem_stage_inst_dmem_n5472,
         mem_stage_inst_dmem_n5471, mem_stage_inst_dmem_n5470,
         mem_stage_inst_dmem_n5469, mem_stage_inst_dmem_n5468,
         mem_stage_inst_dmem_n5467, mem_stage_inst_dmem_n5466,
         mem_stage_inst_dmem_n5465, mem_stage_inst_dmem_n5464,
         mem_stage_inst_dmem_n5463, mem_stage_inst_dmem_n5462,
         mem_stage_inst_dmem_n5461, mem_stage_inst_dmem_n5460,
         mem_stage_inst_dmem_n5459, mem_stage_inst_dmem_n5458,
         mem_stage_inst_dmem_n5457, mem_stage_inst_dmem_n5456,
         mem_stage_inst_dmem_n5455, mem_stage_inst_dmem_n5454,
         mem_stage_inst_dmem_n5453, mem_stage_inst_dmem_n5452,
         mem_stage_inst_dmem_n5451, mem_stage_inst_dmem_n5450,
         mem_stage_inst_dmem_n5449, mem_stage_inst_dmem_n5448,
         mem_stage_inst_dmem_n5447, mem_stage_inst_dmem_n5446,
         mem_stage_inst_dmem_n5445, mem_stage_inst_dmem_n5444,
         mem_stage_inst_dmem_n5443, mem_stage_inst_dmem_n5442,
         mem_stage_inst_dmem_n5441, mem_stage_inst_dmem_n5440,
         mem_stage_inst_dmem_n5439, mem_stage_inst_dmem_n5438,
         mem_stage_inst_dmem_n5437, mem_stage_inst_dmem_n5436,
         mem_stage_inst_dmem_n5435, mem_stage_inst_dmem_n5434,
         mem_stage_inst_dmem_n5433, mem_stage_inst_dmem_n5432,
         mem_stage_inst_dmem_n5431, mem_stage_inst_dmem_n5430,
         mem_stage_inst_dmem_n5429, mem_stage_inst_dmem_n5428,
         mem_stage_inst_dmem_n5427, mem_stage_inst_dmem_n5426,
         mem_stage_inst_dmem_n5425, mem_stage_inst_dmem_n5424,
         mem_stage_inst_dmem_n5423, mem_stage_inst_dmem_n5422,
         mem_stage_inst_dmem_n5421, mem_stage_inst_dmem_n5420,
         mem_stage_inst_dmem_n5419, mem_stage_inst_dmem_n5418,
         mem_stage_inst_dmem_n5417, mem_stage_inst_dmem_n5416,
         mem_stage_inst_dmem_n5415, mem_stage_inst_dmem_n5414,
         mem_stage_inst_dmem_n5413, mem_stage_inst_dmem_n5412,
         mem_stage_inst_dmem_n5411, mem_stage_inst_dmem_n5410,
         mem_stage_inst_dmem_n5409, mem_stage_inst_dmem_n5408,
         mem_stage_inst_dmem_n5407, mem_stage_inst_dmem_n5406,
         mem_stage_inst_dmem_n5405, mem_stage_inst_dmem_n5404,
         mem_stage_inst_dmem_n5403, mem_stage_inst_dmem_n5402,
         mem_stage_inst_dmem_n5401, mem_stage_inst_dmem_n5400,
         mem_stage_inst_dmem_n5399, mem_stage_inst_dmem_n5398,
         mem_stage_inst_dmem_n5397, mem_stage_inst_dmem_n5396,
         mem_stage_inst_dmem_n5395, mem_stage_inst_dmem_n5394,
         mem_stage_inst_dmem_n5393, mem_stage_inst_dmem_n5392,
         mem_stage_inst_dmem_n5391, mem_stage_inst_dmem_n5390,
         mem_stage_inst_dmem_n5389, mem_stage_inst_dmem_n5388,
         mem_stage_inst_dmem_n5387, mem_stage_inst_dmem_n5386,
         mem_stage_inst_dmem_n5385, mem_stage_inst_dmem_n5384,
         mem_stage_inst_dmem_n5383, mem_stage_inst_dmem_n5382,
         mem_stage_inst_dmem_n5381, mem_stage_inst_dmem_n5380,
         mem_stage_inst_dmem_n5379, mem_stage_inst_dmem_n5378,
         mem_stage_inst_dmem_n5377, mem_stage_inst_dmem_n5376,
         mem_stage_inst_dmem_n5375, mem_stage_inst_dmem_n5374,
         mem_stage_inst_dmem_n5373, mem_stage_inst_dmem_n5372,
         mem_stage_inst_dmem_n5371, mem_stage_inst_dmem_n5370,
         mem_stage_inst_dmem_n5369, mem_stage_inst_dmem_n5368,
         mem_stage_inst_dmem_n5367, mem_stage_inst_dmem_n5366,
         mem_stage_inst_dmem_n5365, mem_stage_inst_dmem_n5364,
         mem_stage_inst_dmem_n5363, mem_stage_inst_dmem_n5362,
         mem_stage_inst_dmem_n5361, mem_stage_inst_dmem_n5360,
         mem_stage_inst_dmem_n5359, mem_stage_inst_dmem_n5358,
         mem_stage_inst_dmem_n5357, mem_stage_inst_dmem_n5356,
         mem_stage_inst_dmem_n5355, mem_stage_inst_dmem_n5354,
         mem_stage_inst_dmem_n5353, mem_stage_inst_dmem_n5352,
         mem_stage_inst_dmem_n5351, mem_stage_inst_dmem_n5350,
         mem_stage_inst_dmem_n5349, mem_stage_inst_dmem_n5348,
         mem_stage_inst_dmem_n5347, mem_stage_inst_dmem_n5346,
         mem_stage_inst_dmem_n5345, mem_stage_inst_dmem_n5344,
         mem_stage_inst_dmem_n5343, mem_stage_inst_dmem_n5342,
         mem_stage_inst_dmem_n5341, mem_stage_inst_dmem_n5340,
         mem_stage_inst_dmem_n5339, mem_stage_inst_dmem_n5338,
         mem_stage_inst_dmem_n5337, mem_stage_inst_dmem_n5336,
         mem_stage_inst_dmem_n5335, mem_stage_inst_dmem_n5334,
         mem_stage_inst_dmem_n5333, mem_stage_inst_dmem_n5332,
         mem_stage_inst_dmem_n5331, mem_stage_inst_dmem_n5330,
         mem_stage_inst_dmem_n5329, mem_stage_inst_dmem_n5328,
         mem_stage_inst_dmem_n5327, mem_stage_inst_dmem_n5326,
         mem_stage_inst_dmem_n5325, mem_stage_inst_dmem_n5324,
         mem_stage_inst_dmem_n5323, mem_stage_inst_dmem_n5322,
         mem_stage_inst_dmem_n5321, mem_stage_inst_dmem_n5320,
         mem_stage_inst_dmem_n5319, mem_stage_inst_dmem_n5318,
         mem_stage_inst_dmem_n5317, mem_stage_inst_dmem_n5316,
         mem_stage_inst_dmem_n5315, mem_stage_inst_dmem_n5314,
         mem_stage_inst_dmem_n5313, mem_stage_inst_dmem_n5312,
         mem_stage_inst_dmem_n5311, mem_stage_inst_dmem_n5310,
         mem_stage_inst_dmem_n5309, mem_stage_inst_dmem_n5308,
         mem_stage_inst_dmem_n5307, mem_stage_inst_dmem_n5306,
         mem_stage_inst_dmem_n5305, mem_stage_inst_dmem_n5304,
         mem_stage_inst_dmem_n5303, mem_stage_inst_dmem_n5302,
         mem_stage_inst_dmem_n5301, mem_stage_inst_dmem_n5300,
         mem_stage_inst_dmem_n5299, mem_stage_inst_dmem_n5298,
         mem_stage_inst_dmem_n5297, mem_stage_inst_dmem_n5296,
         mem_stage_inst_dmem_n5295, mem_stage_inst_dmem_n5294,
         mem_stage_inst_dmem_n5293, mem_stage_inst_dmem_n5292,
         mem_stage_inst_dmem_n5291, mem_stage_inst_dmem_n5290,
         mem_stage_inst_dmem_n5289, mem_stage_inst_dmem_n5288,
         mem_stage_inst_dmem_n5287, mem_stage_inst_dmem_n5286,
         mem_stage_inst_dmem_n5285, mem_stage_inst_dmem_n5284,
         mem_stage_inst_dmem_n5283, mem_stage_inst_dmem_n5282,
         mem_stage_inst_dmem_n5281, mem_stage_inst_dmem_n5280,
         mem_stage_inst_dmem_n5279, mem_stage_inst_dmem_n5278,
         mem_stage_inst_dmem_n5277, mem_stage_inst_dmem_n5276,
         mem_stage_inst_dmem_n5275, mem_stage_inst_dmem_n5274,
         mem_stage_inst_dmem_n5273, mem_stage_inst_dmem_n5272,
         mem_stage_inst_dmem_n5271, mem_stage_inst_dmem_n5270,
         mem_stage_inst_dmem_n5269, mem_stage_inst_dmem_n5268,
         mem_stage_inst_dmem_n5267, mem_stage_inst_dmem_n5266,
         mem_stage_inst_dmem_n5265, mem_stage_inst_dmem_n5264,
         mem_stage_inst_dmem_n5263, mem_stage_inst_dmem_n5262,
         mem_stage_inst_dmem_n5261, mem_stage_inst_dmem_n5260,
         mem_stage_inst_dmem_n5259, mem_stage_inst_dmem_n5258,
         mem_stage_inst_dmem_n5257, mem_stage_inst_dmem_n5256,
         mem_stage_inst_dmem_n5255, mem_stage_inst_dmem_n5254,
         mem_stage_inst_dmem_n5253, mem_stage_inst_dmem_n5252,
         mem_stage_inst_dmem_n5251, mem_stage_inst_dmem_n5250,
         mem_stage_inst_dmem_n5249, mem_stage_inst_dmem_n5248,
         mem_stage_inst_dmem_n5247, mem_stage_inst_dmem_n5246,
         mem_stage_inst_dmem_n5245, mem_stage_inst_dmem_n5244,
         mem_stage_inst_dmem_n5243, mem_stage_inst_dmem_n5242,
         mem_stage_inst_dmem_n5241, mem_stage_inst_dmem_n5240,
         mem_stage_inst_dmem_n5239, mem_stage_inst_dmem_n5238,
         mem_stage_inst_dmem_n5237, mem_stage_inst_dmem_n5236,
         mem_stage_inst_dmem_n5235, mem_stage_inst_dmem_n5234,
         mem_stage_inst_dmem_n5233, mem_stage_inst_dmem_n5232,
         mem_stage_inst_dmem_n5231, mem_stage_inst_dmem_n5230,
         mem_stage_inst_dmem_n5229, mem_stage_inst_dmem_n5228,
         mem_stage_inst_dmem_n5227, mem_stage_inst_dmem_n5226,
         mem_stage_inst_dmem_n5225, mem_stage_inst_dmem_n5224,
         mem_stage_inst_dmem_n5223, mem_stage_inst_dmem_n5222,
         mem_stage_inst_dmem_n5221, mem_stage_inst_dmem_n5220,
         mem_stage_inst_dmem_n5219, mem_stage_inst_dmem_n5218,
         mem_stage_inst_dmem_n5217, mem_stage_inst_dmem_n5216,
         mem_stage_inst_dmem_n5215, mem_stage_inst_dmem_n5214,
         mem_stage_inst_dmem_n5213, mem_stage_inst_dmem_n5212,
         mem_stage_inst_dmem_n5211, mem_stage_inst_dmem_n5210,
         mem_stage_inst_dmem_n5209, mem_stage_inst_dmem_n5208,
         mem_stage_inst_dmem_n5207, mem_stage_inst_dmem_n5206,
         mem_stage_inst_dmem_n5205, mem_stage_inst_dmem_n5204,
         mem_stage_inst_dmem_n5203, mem_stage_inst_dmem_n5202,
         mem_stage_inst_dmem_n5201, mem_stage_inst_dmem_n5200,
         mem_stage_inst_dmem_n5199, mem_stage_inst_dmem_n5198,
         mem_stage_inst_dmem_n5197, mem_stage_inst_dmem_n5196,
         mem_stage_inst_dmem_n5195, mem_stage_inst_dmem_n5194,
         mem_stage_inst_dmem_n5193, mem_stage_inst_dmem_n5192,
         mem_stage_inst_dmem_n5191, mem_stage_inst_dmem_n5190,
         mem_stage_inst_dmem_n5189, mem_stage_inst_dmem_n5188,
         mem_stage_inst_dmem_n5187, mem_stage_inst_dmem_n5186,
         mem_stage_inst_dmem_n5185, mem_stage_inst_dmem_n5184,
         mem_stage_inst_dmem_n5183, mem_stage_inst_dmem_n5182,
         mem_stage_inst_dmem_n5181, mem_stage_inst_dmem_n5180,
         mem_stage_inst_dmem_n5179, mem_stage_inst_dmem_n5178,
         mem_stage_inst_dmem_n5177, mem_stage_inst_dmem_n5176,
         mem_stage_inst_dmem_n5175, mem_stage_inst_dmem_n5174,
         mem_stage_inst_dmem_n5173, mem_stage_inst_dmem_n5172,
         mem_stage_inst_dmem_n5171, mem_stage_inst_dmem_n5170,
         mem_stage_inst_dmem_n5169, mem_stage_inst_dmem_n5168,
         mem_stage_inst_dmem_n5167, mem_stage_inst_dmem_n5166,
         mem_stage_inst_dmem_n5165, mem_stage_inst_dmem_n5164,
         mem_stage_inst_dmem_n5163, mem_stage_inst_dmem_n5162,
         mem_stage_inst_dmem_n5161, mem_stage_inst_dmem_n5160,
         mem_stage_inst_dmem_n5159, mem_stage_inst_dmem_n5158,
         mem_stage_inst_dmem_n5157, mem_stage_inst_dmem_n5156,
         mem_stage_inst_dmem_n5155, mem_stage_inst_dmem_n5154,
         mem_stage_inst_dmem_n5153, mem_stage_inst_dmem_n5152,
         mem_stage_inst_dmem_n5151, mem_stage_inst_dmem_n5150,
         mem_stage_inst_dmem_n5149, mem_stage_inst_dmem_n5148,
         mem_stage_inst_dmem_n5147, mem_stage_inst_dmem_n5146,
         mem_stage_inst_dmem_n5145, mem_stage_inst_dmem_n5144,
         mem_stage_inst_dmem_n5143, mem_stage_inst_dmem_n5142,
         mem_stage_inst_dmem_n5141, mem_stage_inst_dmem_n5140,
         mem_stage_inst_dmem_n5139, mem_stage_inst_dmem_n5138,
         mem_stage_inst_dmem_n5137, mem_stage_inst_dmem_n5136,
         mem_stage_inst_dmem_n5135, mem_stage_inst_dmem_n5134,
         mem_stage_inst_dmem_n5133, mem_stage_inst_dmem_n5132,
         mem_stage_inst_dmem_n5131, mem_stage_inst_dmem_n5130,
         mem_stage_inst_dmem_n5129, mem_stage_inst_dmem_n5128,
         mem_stage_inst_dmem_n5127, mem_stage_inst_dmem_n5126,
         mem_stage_inst_dmem_n5125, mem_stage_inst_dmem_n5124,
         mem_stage_inst_dmem_n5123, mem_stage_inst_dmem_n5122,
         mem_stage_inst_dmem_n5121, mem_stage_inst_dmem_n5120,
         mem_stage_inst_dmem_n5119, mem_stage_inst_dmem_n5118,
         mem_stage_inst_dmem_n5117, mem_stage_inst_dmem_n5116,
         mem_stage_inst_dmem_n5115, mem_stage_inst_dmem_n5114,
         mem_stage_inst_dmem_n5113, mem_stage_inst_dmem_n5112,
         mem_stage_inst_dmem_n5111, mem_stage_inst_dmem_n5110,
         mem_stage_inst_dmem_n5109, mem_stage_inst_dmem_n5108,
         mem_stage_inst_dmem_n5107, mem_stage_inst_dmem_n5106,
         mem_stage_inst_dmem_n5105, mem_stage_inst_dmem_n5104,
         mem_stage_inst_dmem_n5103, mem_stage_inst_dmem_n5102,
         mem_stage_inst_dmem_n5101, mem_stage_inst_dmem_n5100,
         mem_stage_inst_dmem_n5099, mem_stage_inst_dmem_n5098,
         mem_stage_inst_dmem_n5097, mem_stage_inst_dmem_n5096,
         mem_stage_inst_dmem_n5095, mem_stage_inst_dmem_n5094,
         mem_stage_inst_dmem_n5093, mem_stage_inst_dmem_n5092,
         mem_stage_inst_dmem_n5091, mem_stage_inst_dmem_n5090,
         mem_stage_inst_dmem_n5089, mem_stage_inst_dmem_n5088,
         mem_stage_inst_dmem_n5087, mem_stage_inst_dmem_n5086,
         mem_stage_inst_dmem_n5085, mem_stage_inst_dmem_n5084,
         mem_stage_inst_dmem_n5083, mem_stage_inst_dmem_n5082,
         mem_stage_inst_dmem_n5081, mem_stage_inst_dmem_n5080,
         mem_stage_inst_dmem_n5079, mem_stage_inst_dmem_n5078,
         mem_stage_inst_dmem_n5077, mem_stage_inst_dmem_n5076,
         mem_stage_inst_dmem_n5075, mem_stage_inst_dmem_n5074,
         mem_stage_inst_dmem_n5073, mem_stage_inst_dmem_n5072,
         mem_stage_inst_dmem_n5071, mem_stage_inst_dmem_n5070,
         mem_stage_inst_dmem_n5069, mem_stage_inst_dmem_n5068,
         mem_stage_inst_dmem_n5067, mem_stage_inst_dmem_n5066,
         mem_stage_inst_dmem_n5065, mem_stage_inst_dmem_n5064,
         mem_stage_inst_dmem_n5063, mem_stage_inst_dmem_n5062,
         mem_stage_inst_dmem_n5061, mem_stage_inst_dmem_n5060,
         mem_stage_inst_dmem_n5059, mem_stage_inst_dmem_n5058,
         mem_stage_inst_dmem_n5057, mem_stage_inst_dmem_n5056,
         mem_stage_inst_dmem_n5055, mem_stage_inst_dmem_n5054,
         mem_stage_inst_dmem_n5053, mem_stage_inst_dmem_n5052,
         mem_stage_inst_dmem_n5051, mem_stage_inst_dmem_n5050,
         mem_stage_inst_dmem_n5049, mem_stage_inst_dmem_n5048,
         mem_stage_inst_dmem_n5047, mem_stage_inst_dmem_n5046,
         mem_stage_inst_dmem_n5045, mem_stage_inst_dmem_n5044,
         mem_stage_inst_dmem_n5043, mem_stage_inst_dmem_n5042,
         mem_stage_inst_dmem_n5041, mem_stage_inst_dmem_n5040,
         mem_stage_inst_dmem_n5039, mem_stage_inst_dmem_n5038,
         mem_stage_inst_dmem_n5037, mem_stage_inst_dmem_n5036,
         mem_stage_inst_dmem_n5035, mem_stage_inst_dmem_n5034,
         mem_stage_inst_dmem_n5033, mem_stage_inst_dmem_n5032,
         mem_stage_inst_dmem_n5031, mem_stage_inst_dmem_n5030,
         mem_stage_inst_dmem_n5029, mem_stage_inst_dmem_n5028,
         mem_stage_inst_dmem_n5027, mem_stage_inst_dmem_n5026,
         mem_stage_inst_dmem_n5025, mem_stage_inst_dmem_n5024,
         mem_stage_inst_dmem_n5023, mem_stage_inst_dmem_n5022,
         mem_stage_inst_dmem_n5021, mem_stage_inst_dmem_n5020,
         mem_stage_inst_dmem_n5019, mem_stage_inst_dmem_n5018,
         mem_stage_inst_dmem_n5017, mem_stage_inst_dmem_n5016,
         mem_stage_inst_dmem_n5015, mem_stage_inst_dmem_n5014,
         mem_stage_inst_dmem_n5013, mem_stage_inst_dmem_n5012,
         mem_stage_inst_dmem_n5011, mem_stage_inst_dmem_n5010,
         mem_stage_inst_dmem_n5009, mem_stage_inst_dmem_n5008,
         mem_stage_inst_dmem_n5007, mem_stage_inst_dmem_n5006,
         mem_stage_inst_dmem_n5005, mem_stage_inst_dmem_n5004,
         mem_stage_inst_dmem_n5003, mem_stage_inst_dmem_n5002,
         mem_stage_inst_dmem_n5001, mem_stage_inst_dmem_n5000,
         mem_stage_inst_dmem_n4999, mem_stage_inst_dmem_n4998,
         mem_stage_inst_dmem_n4997, mem_stage_inst_dmem_n4996,
         mem_stage_inst_dmem_n4995, mem_stage_inst_dmem_n4994,
         mem_stage_inst_dmem_n4993, mem_stage_inst_dmem_n4992,
         mem_stage_inst_dmem_n4991, mem_stage_inst_dmem_n4990,
         mem_stage_inst_dmem_n4989, mem_stage_inst_dmem_n4988,
         mem_stage_inst_dmem_n4987, mem_stage_inst_dmem_n4986,
         mem_stage_inst_dmem_n4985, mem_stage_inst_dmem_n4984,
         mem_stage_inst_dmem_n4983, mem_stage_inst_dmem_n4982,
         mem_stage_inst_dmem_n4981, mem_stage_inst_dmem_n4980,
         mem_stage_inst_dmem_n4979, mem_stage_inst_dmem_n4978,
         mem_stage_inst_dmem_n4977, mem_stage_inst_dmem_n4976,
         mem_stage_inst_dmem_n4975, mem_stage_inst_dmem_n4974,
         mem_stage_inst_dmem_n4973, mem_stage_inst_dmem_n4972,
         mem_stage_inst_dmem_n4971, mem_stage_inst_dmem_n4970,
         mem_stage_inst_dmem_n4969, mem_stage_inst_dmem_n4968,
         mem_stage_inst_dmem_n4967, mem_stage_inst_dmem_n4966,
         mem_stage_inst_dmem_n4965, mem_stage_inst_dmem_n4964,
         mem_stage_inst_dmem_n4963, mem_stage_inst_dmem_n4962,
         mem_stage_inst_dmem_n4961, mem_stage_inst_dmem_n4960,
         mem_stage_inst_dmem_n4959, mem_stage_inst_dmem_n4958,
         mem_stage_inst_dmem_n4957, mem_stage_inst_dmem_n4956,
         mem_stage_inst_dmem_n4955, mem_stage_inst_dmem_n4954,
         mem_stage_inst_dmem_n4953, mem_stage_inst_dmem_n4952,
         mem_stage_inst_dmem_n4951, mem_stage_inst_dmem_n4950,
         mem_stage_inst_dmem_n4949, mem_stage_inst_dmem_n4948,
         mem_stage_inst_dmem_n4947, mem_stage_inst_dmem_n4946,
         mem_stage_inst_dmem_n4945, mem_stage_inst_dmem_n4944,
         mem_stage_inst_dmem_n4943, mem_stage_inst_dmem_n4942,
         mem_stage_inst_dmem_n4941, mem_stage_inst_dmem_n4940,
         mem_stage_inst_dmem_n4939, mem_stage_inst_dmem_n4938,
         mem_stage_inst_dmem_n4937, mem_stage_inst_dmem_n4936,
         mem_stage_inst_dmem_n4935, mem_stage_inst_dmem_n4934,
         mem_stage_inst_dmem_n4933, mem_stage_inst_dmem_n4932,
         mem_stage_inst_dmem_n4931, mem_stage_inst_dmem_n4930,
         mem_stage_inst_dmem_n4929, mem_stage_inst_dmem_n4928,
         mem_stage_inst_dmem_n4927, mem_stage_inst_dmem_n4926,
         mem_stage_inst_dmem_n4925, mem_stage_inst_dmem_n4924,
         mem_stage_inst_dmem_n4923, mem_stage_inst_dmem_n4922,
         mem_stage_inst_dmem_n4921, mem_stage_inst_dmem_n4920,
         mem_stage_inst_dmem_n4919, mem_stage_inst_dmem_n4918,
         mem_stage_inst_dmem_n4917, mem_stage_inst_dmem_n4916,
         mem_stage_inst_dmem_n4915, mem_stage_inst_dmem_n4914,
         mem_stage_inst_dmem_n4913, mem_stage_inst_dmem_n4912,
         mem_stage_inst_dmem_n4911, mem_stage_inst_dmem_n4910,
         mem_stage_inst_dmem_n4909, mem_stage_inst_dmem_n4908,
         mem_stage_inst_dmem_n4907, mem_stage_inst_dmem_n4906,
         mem_stage_inst_dmem_n4905, mem_stage_inst_dmem_n4904,
         mem_stage_inst_dmem_n4903, mem_stage_inst_dmem_n4902,
         mem_stage_inst_dmem_n4901, mem_stage_inst_dmem_n4900,
         mem_stage_inst_dmem_n4899, mem_stage_inst_dmem_n4898,
         mem_stage_inst_dmem_n4897, mem_stage_inst_dmem_n4896,
         mem_stage_inst_dmem_n4895, mem_stage_inst_dmem_n4894,
         mem_stage_inst_dmem_n4893, mem_stage_inst_dmem_n4892,
         mem_stage_inst_dmem_n4891, mem_stage_inst_dmem_n4890,
         mem_stage_inst_dmem_n4889, mem_stage_inst_dmem_n4888,
         mem_stage_inst_dmem_n4887, mem_stage_inst_dmem_n4886,
         mem_stage_inst_dmem_n4885, mem_stage_inst_dmem_n4884,
         mem_stage_inst_dmem_n4883, mem_stage_inst_dmem_n4882,
         mem_stage_inst_dmem_n4881, mem_stage_inst_dmem_n4880,
         mem_stage_inst_dmem_n4879, mem_stage_inst_dmem_n4878,
         mem_stage_inst_dmem_n4877, mem_stage_inst_dmem_n4876,
         mem_stage_inst_dmem_n4875, mem_stage_inst_dmem_n4874,
         mem_stage_inst_dmem_n4873, mem_stage_inst_dmem_n4872,
         mem_stage_inst_dmem_n4871, mem_stage_inst_dmem_n4870,
         mem_stage_inst_dmem_n4869, mem_stage_inst_dmem_n4868,
         mem_stage_inst_dmem_n4867, mem_stage_inst_dmem_n4866,
         mem_stage_inst_dmem_n4865, mem_stage_inst_dmem_n4864,
         mem_stage_inst_dmem_n4863, mem_stage_inst_dmem_n4862,
         mem_stage_inst_dmem_n4861, mem_stage_inst_dmem_n4860,
         mem_stage_inst_dmem_n4859, mem_stage_inst_dmem_n4858,
         mem_stage_inst_dmem_n4857, mem_stage_inst_dmem_n4856,
         mem_stage_inst_dmem_n4855, mem_stage_inst_dmem_n4854,
         mem_stage_inst_dmem_n4853, mem_stage_inst_dmem_n4852,
         mem_stage_inst_dmem_n4851, mem_stage_inst_dmem_n4850,
         mem_stage_inst_dmem_n4849, mem_stage_inst_dmem_n4848,
         mem_stage_inst_dmem_n4847, mem_stage_inst_dmem_n4846,
         mem_stage_inst_dmem_n4845, mem_stage_inst_dmem_n4844,
         mem_stage_inst_dmem_n4843, mem_stage_inst_dmem_n4842,
         mem_stage_inst_dmem_n4841, mem_stage_inst_dmem_n4840,
         mem_stage_inst_dmem_n4839, mem_stage_inst_dmem_n4838,
         mem_stage_inst_dmem_n4837, mem_stage_inst_dmem_n4836,
         mem_stage_inst_dmem_n4835, mem_stage_inst_dmem_n4834,
         mem_stage_inst_dmem_n4833, mem_stage_inst_dmem_n4832,
         mem_stage_inst_dmem_n4831, mem_stage_inst_dmem_n4830,
         mem_stage_inst_dmem_n4829, mem_stage_inst_dmem_n4828,
         mem_stage_inst_dmem_n4827, mem_stage_inst_dmem_n4826,
         mem_stage_inst_dmem_n4825, mem_stage_inst_dmem_n4824,
         mem_stage_inst_dmem_n4823, mem_stage_inst_dmem_n4822,
         mem_stage_inst_dmem_n4821, mem_stage_inst_dmem_n4820,
         mem_stage_inst_dmem_n4819, mem_stage_inst_dmem_n4818,
         mem_stage_inst_dmem_n4817, mem_stage_inst_dmem_n4816,
         mem_stage_inst_dmem_n4815, mem_stage_inst_dmem_n4814,
         mem_stage_inst_dmem_n4813, mem_stage_inst_dmem_n4812,
         mem_stage_inst_dmem_n4811, mem_stage_inst_dmem_n4810,
         mem_stage_inst_dmem_n4809, mem_stage_inst_dmem_n4808,
         mem_stage_inst_dmem_n4807, mem_stage_inst_dmem_n4806,
         mem_stage_inst_dmem_n4805, mem_stage_inst_dmem_n4804,
         mem_stage_inst_dmem_n4803, mem_stage_inst_dmem_n4802,
         mem_stage_inst_dmem_n4801, mem_stage_inst_dmem_n4800,
         mem_stage_inst_dmem_n4799, mem_stage_inst_dmem_n4798,
         mem_stage_inst_dmem_n4797, mem_stage_inst_dmem_n4796,
         mem_stage_inst_dmem_n4795, mem_stage_inst_dmem_n4794,
         mem_stage_inst_dmem_n4793, mem_stage_inst_dmem_n4792,
         mem_stage_inst_dmem_n4791, mem_stage_inst_dmem_n4790,
         mem_stage_inst_dmem_n4789, mem_stage_inst_dmem_n4788,
         mem_stage_inst_dmem_n4787, mem_stage_inst_dmem_n4786,
         mem_stage_inst_dmem_n4785, mem_stage_inst_dmem_n4784,
         mem_stage_inst_dmem_n4783, mem_stage_inst_dmem_n4782,
         mem_stage_inst_dmem_n4781, mem_stage_inst_dmem_n4780,
         mem_stage_inst_dmem_n4779, mem_stage_inst_dmem_n4778,
         mem_stage_inst_dmem_n4777, mem_stage_inst_dmem_n4776,
         mem_stage_inst_dmem_n4775, mem_stage_inst_dmem_n4774,
         mem_stage_inst_dmem_n4773, mem_stage_inst_dmem_n4772,
         mem_stage_inst_dmem_n4771, mem_stage_inst_dmem_n4770,
         mem_stage_inst_dmem_n4769, mem_stage_inst_dmem_n4768,
         mem_stage_inst_dmem_n4767, mem_stage_inst_dmem_n4766,
         mem_stage_inst_dmem_n4765, mem_stage_inst_dmem_n4764,
         mem_stage_inst_dmem_n4763, mem_stage_inst_dmem_n4762,
         mem_stage_inst_dmem_n4761, mem_stage_inst_dmem_n4760,
         mem_stage_inst_dmem_n4759, mem_stage_inst_dmem_n4758,
         mem_stage_inst_dmem_n4757, mem_stage_inst_dmem_n4756,
         mem_stage_inst_dmem_n4755, mem_stage_inst_dmem_n4754,
         mem_stage_inst_dmem_n4753, mem_stage_inst_dmem_n4752,
         mem_stage_inst_dmem_n4751, mem_stage_inst_dmem_n4750,
         mem_stage_inst_dmem_n4749, mem_stage_inst_dmem_n4748,
         mem_stage_inst_dmem_n4747, mem_stage_inst_dmem_n4746,
         mem_stage_inst_dmem_n4745, mem_stage_inst_dmem_n4744,
         mem_stage_inst_dmem_n4743, mem_stage_inst_dmem_n4742,
         mem_stage_inst_dmem_n4741, mem_stage_inst_dmem_n4740,
         mem_stage_inst_dmem_n4739, mem_stage_inst_dmem_n4738,
         mem_stage_inst_dmem_n4737, mem_stage_inst_dmem_n4736,
         mem_stage_inst_dmem_n4735, mem_stage_inst_dmem_n4734,
         mem_stage_inst_dmem_n4733, mem_stage_inst_dmem_n4732,
         mem_stage_inst_dmem_n4731, mem_stage_inst_dmem_n4730,
         mem_stage_inst_dmem_n4729, mem_stage_inst_dmem_n4728,
         mem_stage_inst_dmem_n4727, mem_stage_inst_dmem_n4726,
         mem_stage_inst_dmem_n4725, mem_stage_inst_dmem_n4724,
         mem_stage_inst_dmem_n4723, mem_stage_inst_dmem_n4722,
         mem_stage_inst_dmem_n4721, mem_stage_inst_dmem_n4720,
         mem_stage_inst_dmem_n4719, mem_stage_inst_dmem_n4718,
         mem_stage_inst_dmem_n4717, mem_stage_inst_dmem_n4716,
         mem_stage_inst_dmem_n4715, mem_stage_inst_dmem_n4714,
         mem_stage_inst_dmem_n4713, mem_stage_inst_dmem_n4712,
         mem_stage_inst_dmem_n4711, mem_stage_inst_dmem_n4710,
         mem_stage_inst_dmem_n4709, mem_stage_inst_dmem_n4708,
         mem_stage_inst_dmem_n4707, mem_stage_inst_dmem_n4706,
         mem_stage_inst_dmem_n4705, mem_stage_inst_dmem_n4704,
         mem_stage_inst_dmem_n4703, mem_stage_inst_dmem_n4702,
         mem_stage_inst_dmem_n4701, mem_stage_inst_dmem_n4700,
         mem_stage_inst_dmem_n4699, mem_stage_inst_dmem_n4698,
         mem_stage_inst_dmem_n4697, mem_stage_inst_dmem_n4696,
         mem_stage_inst_dmem_n4695, mem_stage_inst_dmem_n4694,
         mem_stage_inst_dmem_n4693, mem_stage_inst_dmem_n4692,
         mem_stage_inst_dmem_n4691, mem_stage_inst_dmem_n4690,
         mem_stage_inst_dmem_n4689, mem_stage_inst_dmem_n4688,
         mem_stage_inst_dmem_n4687, mem_stage_inst_dmem_n4686,
         mem_stage_inst_dmem_n4685, mem_stage_inst_dmem_n4684,
         mem_stage_inst_dmem_n4683, mem_stage_inst_dmem_n4682,
         mem_stage_inst_dmem_n4681, mem_stage_inst_dmem_n4680,
         mem_stage_inst_dmem_n4679, mem_stage_inst_dmem_n4678,
         mem_stage_inst_dmem_n4677, mem_stage_inst_dmem_n4676,
         mem_stage_inst_dmem_n4675, mem_stage_inst_dmem_n4674,
         mem_stage_inst_dmem_n4673, mem_stage_inst_dmem_n4672,
         mem_stage_inst_dmem_n4671, mem_stage_inst_dmem_n4670,
         mem_stage_inst_dmem_n4669, mem_stage_inst_dmem_n4668,
         mem_stage_inst_dmem_n4667, mem_stage_inst_dmem_n4666,
         mem_stage_inst_dmem_n4665, mem_stage_inst_dmem_n4664,
         mem_stage_inst_dmem_n4663, mem_stage_inst_dmem_n4662,
         mem_stage_inst_dmem_n4661, mem_stage_inst_dmem_n564,
         mem_stage_inst_dmem_n563, mem_stage_inst_dmem_n562,
         mem_stage_inst_dmem_n561, mem_stage_inst_dmem_n560,
         mem_stage_inst_dmem_n559, mem_stage_inst_dmem_n558,
         mem_stage_inst_dmem_n557, mem_stage_inst_dmem_n556,
         mem_stage_inst_dmem_n555, mem_stage_inst_dmem_n554,
         mem_stage_inst_dmem_n553, mem_stage_inst_dmem_n552,
         mem_stage_inst_dmem_n551, mem_stage_inst_dmem_n550,
         mem_stage_inst_dmem_n549, mem_stage_inst_dmem_n548,
         mem_stage_inst_dmem_n547, mem_stage_inst_dmem_n546,
         mem_stage_inst_dmem_n545, mem_stage_inst_dmem_n544,
         mem_stage_inst_dmem_n543, mem_stage_inst_dmem_n542,
         mem_stage_inst_dmem_n541, mem_stage_inst_dmem_n540,
         mem_stage_inst_dmem_n539, mem_stage_inst_dmem_n538,
         mem_stage_inst_dmem_n537, mem_stage_inst_dmem_n536,
         mem_stage_inst_dmem_n535, mem_stage_inst_dmem_n534,
         mem_stage_inst_dmem_n533, mem_stage_inst_dmem_n532,
         mem_stage_inst_dmem_n531, mem_stage_inst_dmem_n530,
         mem_stage_inst_dmem_n529, mem_stage_inst_dmem_n528,
         mem_stage_inst_dmem_n527, mem_stage_inst_dmem_n526,
         mem_stage_inst_dmem_n525, mem_stage_inst_dmem_n524,
         mem_stage_inst_dmem_n523, mem_stage_inst_dmem_n522,
         mem_stage_inst_dmem_n521, mem_stage_inst_dmem_n520,
         mem_stage_inst_dmem_n519, mem_stage_inst_dmem_n518,
         mem_stage_inst_dmem_n517, mem_stage_inst_dmem_n516,
         mem_stage_inst_dmem_n515, mem_stage_inst_dmem_n514,
         mem_stage_inst_dmem_n513, mem_stage_inst_dmem_n512,
         mem_stage_inst_dmem_n511, mem_stage_inst_dmem_n510,
         mem_stage_inst_dmem_n509, mem_stage_inst_dmem_n508,
         mem_stage_inst_dmem_n507, mem_stage_inst_dmem_n506,
         mem_stage_inst_dmem_n505, mem_stage_inst_dmem_n504,
         mem_stage_inst_dmem_n503, mem_stage_inst_dmem_n502,
         mem_stage_inst_dmem_n501, mem_stage_inst_dmem_n500,
         mem_stage_inst_dmem_n499, mem_stage_inst_dmem_n498,
         mem_stage_inst_dmem_n497, mem_stage_inst_dmem_n496,
         mem_stage_inst_dmem_n495, mem_stage_inst_dmem_n494,
         mem_stage_inst_dmem_n493, mem_stage_inst_dmem_n492,
         mem_stage_inst_dmem_n491, mem_stage_inst_dmem_n490,
         mem_stage_inst_dmem_n489, mem_stage_inst_dmem_n488,
         mem_stage_inst_dmem_n487, mem_stage_inst_dmem_n486,
         mem_stage_inst_dmem_n485, mem_stage_inst_dmem_n484,
         mem_stage_inst_dmem_n483, mem_stage_inst_dmem_n482,
         mem_stage_inst_dmem_n481, mem_stage_inst_dmem_n480,
         mem_stage_inst_dmem_n479, mem_stage_inst_dmem_n478,
         mem_stage_inst_dmem_n477, mem_stage_inst_dmem_n476,
         mem_stage_inst_dmem_n475, mem_stage_inst_dmem_n474,
         mem_stage_inst_dmem_n473, mem_stage_inst_dmem_n472,
         mem_stage_inst_dmem_n471, mem_stage_inst_dmem_n470,
         mem_stage_inst_dmem_n469, mem_stage_inst_dmem_n468,
         mem_stage_inst_dmem_n467, mem_stage_inst_dmem_n466,
         mem_stage_inst_dmem_n465, mem_stage_inst_dmem_n464,
         mem_stage_inst_dmem_n463, mem_stage_inst_dmem_n462,
         mem_stage_inst_dmem_n461, mem_stage_inst_dmem_n460,
         mem_stage_inst_dmem_n459, mem_stage_inst_dmem_n458,
         mem_stage_inst_dmem_n457, mem_stage_inst_dmem_n456,
         mem_stage_inst_dmem_n455, mem_stage_inst_dmem_n454,
         mem_stage_inst_dmem_n453, mem_stage_inst_dmem_n452,
         mem_stage_inst_dmem_n451, mem_stage_inst_dmem_n450,
         mem_stage_inst_dmem_n449, mem_stage_inst_dmem_n448,
         mem_stage_inst_dmem_n447, mem_stage_inst_dmem_n446,
         mem_stage_inst_dmem_n445, mem_stage_inst_dmem_n444,
         mem_stage_inst_dmem_n443, mem_stage_inst_dmem_n442,
         mem_stage_inst_dmem_n441, mem_stage_inst_dmem_n440,
         mem_stage_inst_dmem_n439, mem_stage_inst_dmem_n438,
         mem_stage_inst_dmem_n437, mem_stage_inst_dmem_n436,
         mem_stage_inst_dmem_n435, mem_stage_inst_dmem_n434,
         mem_stage_inst_dmem_n433, mem_stage_inst_dmem_n432,
         mem_stage_inst_dmem_n431, mem_stage_inst_dmem_n430,
         mem_stage_inst_dmem_n429, mem_stage_inst_dmem_n428,
         mem_stage_inst_dmem_n427, mem_stage_inst_dmem_n426,
         mem_stage_inst_dmem_n425, mem_stage_inst_dmem_n424,
         mem_stage_inst_dmem_n423, mem_stage_inst_dmem_n422,
         mem_stage_inst_dmem_n421, mem_stage_inst_dmem_n420,
         mem_stage_inst_dmem_n419, mem_stage_inst_dmem_n418,
         mem_stage_inst_dmem_n417, mem_stage_inst_dmem_n416,
         mem_stage_inst_dmem_n415, mem_stage_inst_dmem_n414,
         mem_stage_inst_dmem_n413, mem_stage_inst_dmem_n412,
         mem_stage_inst_dmem_n411, mem_stage_inst_dmem_n410,
         mem_stage_inst_dmem_n409, mem_stage_inst_dmem_n408,
         mem_stage_inst_dmem_n407, mem_stage_inst_dmem_n406,
         mem_stage_inst_dmem_n405, mem_stage_inst_dmem_n404,
         mem_stage_inst_dmem_n403, mem_stage_inst_dmem_n402,
         mem_stage_inst_dmem_n401, mem_stage_inst_dmem_n400,
         mem_stage_inst_dmem_n399, mem_stage_inst_dmem_n398,
         mem_stage_inst_dmem_n397, mem_stage_inst_dmem_n396,
         mem_stage_inst_dmem_n395, mem_stage_inst_dmem_n394,
         mem_stage_inst_dmem_n393, mem_stage_inst_dmem_n392,
         mem_stage_inst_dmem_n391, mem_stage_inst_dmem_n390,
         mem_stage_inst_dmem_n389, mem_stage_inst_dmem_n388,
         mem_stage_inst_dmem_n387, mem_stage_inst_dmem_n386,
         mem_stage_inst_dmem_n385, mem_stage_inst_dmem_n384,
         mem_stage_inst_dmem_n383, mem_stage_inst_dmem_n382,
         mem_stage_inst_dmem_n381, mem_stage_inst_dmem_n380,
         mem_stage_inst_dmem_n379, mem_stage_inst_dmem_n378,
         mem_stage_inst_dmem_n377, mem_stage_inst_dmem_n376,
         mem_stage_inst_dmem_n375, mem_stage_inst_dmem_n374,
         mem_stage_inst_dmem_n373, mem_stage_inst_dmem_n372,
         mem_stage_inst_dmem_n371, mem_stage_inst_dmem_n370,
         mem_stage_inst_dmem_n369, mem_stage_inst_dmem_n368,
         mem_stage_inst_dmem_n367, mem_stage_inst_dmem_n366,
         mem_stage_inst_dmem_n365, mem_stage_inst_dmem_n364,
         mem_stage_inst_dmem_n363, mem_stage_inst_dmem_n362,
         mem_stage_inst_dmem_n361, mem_stage_inst_dmem_n360,
         mem_stage_inst_dmem_n359, mem_stage_inst_dmem_n358,
         mem_stage_inst_dmem_n357, mem_stage_inst_dmem_n356,
         mem_stage_inst_dmem_n355, mem_stage_inst_dmem_n354,
         mem_stage_inst_dmem_n353, mem_stage_inst_dmem_n352,
         mem_stage_inst_dmem_n351, mem_stage_inst_dmem_n350,
         mem_stage_inst_dmem_n349, mem_stage_inst_dmem_n348,
         mem_stage_inst_dmem_n347, mem_stage_inst_dmem_n346,
         mem_stage_inst_dmem_n345, mem_stage_inst_dmem_n344,
         mem_stage_inst_dmem_n343, mem_stage_inst_dmem_n342,
         mem_stage_inst_dmem_n341, mem_stage_inst_dmem_n340,
         mem_stage_inst_dmem_n339, mem_stage_inst_dmem_n338,
         mem_stage_inst_dmem_n337, mem_stage_inst_dmem_n336,
         mem_stage_inst_dmem_n335, mem_stage_inst_dmem_n334,
         mem_stage_inst_dmem_n333, mem_stage_inst_dmem_n332,
         mem_stage_inst_dmem_n331, mem_stage_inst_dmem_n330,
         mem_stage_inst_dmem_n329, mem_stage_inst_dmem_n328,
         mem_stage_inst_dmem_n327, mem_stage_inst_dmem_n326,
         mem_stage_inst_dmem_n325, mem_stage_inst_dmem_n324,
         mem_stage_inst_dmem_n323, mem_stage_inst_dmem_n322,
         mem_stage_inst_dmem_n321, mem_stage_inst_dmem_n320,
         mem_stage_inst_dmem_n319, mem_stage_inst_dmem_n318,
         mem_stage_inst_dmem_n317, mem_stage_inst_dmem_n316,
         mem_stage_inst_dmem_n315, mem_stage_inst_dmem_n314,
         mem_stage_inst_dmem_n313, mem_stage_inst_dmem_n312,
         mem_stage_inst_dmem_n311, mem_stage_inst_dmem_n310,
         mem_stage_inst_dmem_n309, mem_stage_inst_dmem_n308,
         mem_stage_inst_dmem_n307, mem_stage_inst_dmem_n306,
         mem_stage_inst_dmem_n305, mem_stage_inst_dmem_n304,
         mem_stage_inst_dmem_n303, mem_stage_inst_dmem_n302,
         mem_stage_inst_dmem_n301, mem_stage_inst_dmem_n300,
         mem_stage_inst_dmem_n299, mem_stage_inst_dmem_n298,
         mem_stage_inst_dmem_n297, mem_stage_inst_dmem_n296,
         mem_stage_inst_dmem_n295, mem_stage_inst_dmem_n294,
         mem_stage_inst_dmem_n293, mem_stage_inst_dmem_n292,
         mem_stage_inst_dmem_n291, mem_stage_inst_dmem_n290,
         mem_stage_inst_dmem_n289, mem_stage_inst_dmem_n288,
         mem_stage_inst_dmem_n287, mem_stage_inst_dmem_n286,
         mem_stage_inst_dmem_n285, mem_stage_inst_dmem_n284,
         mem_stage_inst_dmem_n283, mem_stage_inst_dmem_n282,
         mem_stage_inst_dmem_n281, mem_stage_inst_dmem_n280,
         mem_stage_inst_dmem_n279, mem_stage_inst_dmem_n278,
         mem_stage_inst_dmem_n277, mem_stage_inst_dmem_n276,
         mem_stage_inst_dmem_n275, mem_stage_inst_dmem_n274,
         mem_stage_inst_dmem_n273, mem_stage_inst_dmem_n272,
         mem_stage_inst_dmem_n271, mem_stage_inst_dmem_n270,
         mem_stage_inst_dmem_n269, mem_stage_inst_dmem_n268,
         mem_stage_inst_dmem_n267, mem_stage_inst_dmem_n266,
         mem_stage_inst_dmem_n265, mem_stage_inst_dmem_n264,
         mem_stage_inst_dmem_n263, mem_stage_inst_dmem_n262,
         mem_stage_inst_dmem_n261, mem_stage_inst_dmem_n260,
         mem_stage_inst_dmem_n259, mem_stage_inst_dmem_n258,
         mem_stage_inst_dmem_n257, mem_stage_inst_dmem_n256,
         mem_stage_inst_dmem_n255, mem_stage_inst_dmem_n254,
         mem_stage_inst_dmem_n253, mem_stage_inst_dmem_n252,
         mem_stage_inst_dmem_n251, mem_stage_inst_dmem_n250,
         mem_stage_inst_dmem_n249, mem_stage_inst_dmem_n248,
         mem_stage_inst_dmem_n247, mem_stage_inst_dmem_n246,
         mem_stage_inst_dmem_n245, mem_stage_inst_dmem_n244,
         mem_stage_inst_dmem_n243, mem_stage_inst_dmem_n242,
         mem_stage_inst_dmem_n241, mem_stage_inst_dmem_n240,
         mem_stage_inst_dmem_n239, mem_stage_inst_dmem_n238,
         mem_stage_inst_dmem_n237, mem_stage_inst_dmem_n236,
         mem_stage_inst_dmem_n235, mem_stage_inst_dmem_n234,
         mem_stage_inst_dmem_n233, mem_stage_inst_dmem_n232,
         mem_stage_inst_dmem_n231, mem_stage_inst_dmem_n230,
         mem_stage_inst_dmem_n229, mem_stage_inst_dmem_n228,
         mem_stage_inst_dmem_n227, mem_stage_inst_dmem_n226,
         mem_stage_inst_dmem_n225, mem_stage_inst_dmem_n224,
         mem_stage_inst_dmem_n223, mem_stage_inst_dmem_n222,
         mem_stage_inst_dmem_n221, mem_stage_inst_dmem_n220,
         mem_stage_inst_dmem_n219, mem_stage_inst_dmem_n218,
         mem_stage_inst_dmem_n217, mem_stage_inst_dmem_n216,
         mem_stage_inst_dmem_n215, mem_stage_inst_dmem_n214,
         mem_stage_inst_dmem_n213, mem_stage_inst_dmem_n212,
         mem_stage_inst_dmem_n211, mem_stage_inst_dmem_n210,
         mem_stage_inst_dmem_n209, mem_stage_inst_dmem_n208,
         mem_stage_inst_dmem_n207, mem_stage_inst_dmem_n206,
         mem_stage_inst_dmem_n205, mem_stage_inst_dmem_n204,
         mem_stage_inst_dmem_n203, mem_stage_inst_dmem_n202,
         mem_stage_inst_dmem_n201, mem_stage_inst_dmem_n200,
         mem_stage_inst_dmem_n199, mem_stage_inst_dmem_n198,
         mem_stage_inst_dmem_n197, mem_stage_inst_dmem_n196,
         mem_stage_inst_dmem_n195, mem_stage_inst_dmem_n194,
         mem_stage_inst_dmem_n193, mem_stage_inst_dmem_n192,
         mem_stage_inst_dmem_n191, mem_stage_inst_dmem_n190,
         mem_stage_inst_dmem_n189, mem_stage_inst_dmem_n188,
         mem_stage_inst_dmem_n187, mem_stage_inst_dmem_n186,
         mem_stage_inst_dmem_n185, mem_stage_inst_dmem_n184,
         mem_stage_inst_dmem_n183, mem_stage_inst_dmem_n182,
         mem_stage_inst_dmem_n181, mem_stage_inst_dmem_n180,
         mem_stage_inst_dmem_n179, mem_stage_inst_dmem_n178,
         mem_stage_inst_dmem_n177, mem_stage_inst_dmem_n176,
         mem_stage_inst_dmem_n175, mem_stage_inst_dmem_n174,
         mem_stage_inst_dmem_n173, mem_stage_inst_dmem_n172,
         mem_stage_inst_dmem_n171, mem_stage_inst_dmem_n170,
         mem_stage_inst_dmem_n169, mem_stage_inst_dmem_n168,
         mem_stage_inst_dmem_n167, mem_stage_inst_dmem_n166,
         mem_stage_inst_dmem_n165, mem_stage_inst_dmem_n164,
         mem_stage_inst_dmem_n163, mem_stage_inst_dmem_n162,
         mem_stage_inst_dmem_n161, mem_stage_inst_dmem_n160,
         mem_stage_inst_dmem_n159, mem_stage_inst_dmem_n158,
         mem_stage_inst_dmem_n157, mem_stage_inst_dmem_n156,
         mem_stage_inst_dmem_n155, mem_stage_inst_dmem_n154,
         mem_stage_inst_dmem_n153, mem_stage_inst_dmem_n152,
         mem_stage_inst_dmem_n151, mem_stage_inst_dmem_n150,
         mem_stage_inst_dmem_n149, mem_stage_inst_dmem_n148,
         mem_stage_inst_dmem_n147, mem_stage_inst_dmem_n146,
         mem_stage_inst_dmem_n145, mem_stage_inst_dmem_n144,
         mem_stage_inst_dmem_n143, mem_stage_inst_dmem_n142,
         mem_stage_inst_dmem_n141, mem_stage_inst_dmem_n140,
         mem_stage_inst_dmem_n139, mem_stage_inst_dmem_n138,
         mem_stage_inst_dmem_n137, mem_stage_inst_dmem_n136,
         mem_stage_inst_dmem_n135, mem_stage_inst_dmem_n134,
         mem_stage_inst_dmem_n133, mem_stage_inst_dmem_n132,
         mem_stage_inst_dmem_n131, mem_stage_inst_dmem_n130,
         mem_stage_inst_dmem_n129, mem_stage_inst_dmem_n128,
         mem_stage_inst_dmem_n127, mem_stage_inst_dmem_n126,
         mem_stage_inst_dmem_n125, mem_stage_inst_dmem_n124,
         mem_stage_inst_dmem_n123, mem_stage_inst_dmem_n122,
         mem_stage_inst_dmem_n121, mem_stage_inst_dmem_n120,
         mem_stage_inst_dmem_n119, mem_stage_inst_dmem_n118,
         mem_stage_inst_dmem_n117, mem_stage_inst_dmem_n116,
         mem_stage_inst_dmem_n115, mem_stage_inst_dmem_n114,
         mem_stage_inst_dmem_n113, mem_stage_inst_dmem_n112,
         mem_stage_inst_dmem_n111, mem_stage_inst_dmem_n110,
         mem_stage_inst_dmem_n109, mem_stage_inst_dmem_n108,
         mem_stage_inst_dmem_n107, mem_stage_inst_dmem_n106,
         mem_stage_inst_dmem_n105, mem_stage_inst_dmem_n104,
         mem_stage_inst_dmem_n103, mem_stage_inst_dmem_n102,
         mem_stage_inst_dmem_n101, mem_stage_inst_dmem_n100,
         mem_stage_inst_dmem_n99, mem_stage_inst_dmem_n98,
         mem_stage_inst_dmem_n97, mem_stage_inst_dmem_n96,
         mem_stage_inst_dmem_n95, mem_stage_inst_dmem_n94,
         mem_stage_inst_dmem_n93, mem_stage_inst_dmem_n92,
         mem_stage_inst_dmem_n91, mem_stage_inst_dmem_n90,
         mem_stage_inst_dmem_n89, mem_stage_inst_dmem_n88,
         mem_stage_inst_dmem_n87, mem_stage_inst_dmem_n86,
         mem_stage_inst_dmem_n85, mem_stage_inst_dmem_n84,
         mem_stage_inst_dmem_n83, mem_stage_inst_dmem_n82,
         mem_stage_inst_dmem_n81, mem_stage_inst_dmem_n80,
         mem_stage_inst_dmem_n79, mem_stage_inst_dmem_n78,
         mem_stage_inst_dmem_n77, mem_stage_inst_dmem_n76,
         mem_stage_inst_dmem_n75, mem_stage_inst_dmem_n74,
         mem_stage_inst_dmem_n73, mem_stage_inst_dmem_n72,
         mem_stage_inst_dmem_n71, mem_stage_inst_dmem_n70,
         mem_stage_inst_dmem_n69, mem_stage_inst_dmem_n68,
         mem_stage_inst_dmem_n67, mem_stage_inst_dmem_n66,
         mem_stage_inst_dmem_n65, mem_stage_inst_dmem_n64,
         mem_stage_inst_dmem_n63, mem_stage_inst_dmem_n62,
         mem_stage_inst_dmem_n61, mem_stage_inst_dmem_n60,
         mem_stage_inst_dmem_n59, mem_stage_inst_dmem_n58,
         mem_stage_inst_dmem_n57, mem_stage_inst_dmem_n56,
         mem_stage_inst_dmem_n55, mem_stage_inst_dmem_n54,
         mem_stage_inst_dmem_n53, mem_stage_inst_dmem_n52,
         mem_stage_inst_dmem_n51, mem_stage_inst_dmem_n50,
         mem_stage_inst_dmem_n49, mem_stage_inst_dmem_n48,
         mem_stage_inst_dmem_n47, mem_stage_inst_dmem_n46,
         mem_stage_inst_dmem_n45, mem_stage_inst_dmem_n44,
         mem_stage_inst_dmem_n43, mem_stage_inst_dmem_n42,
         mem_stage_inst_dmem_n41, mem_stage_inst_dmem_n40,
         mem_stage_inst_dmem_n39, mem_stage_inst_dmem_n38,
         mem_stage_inst_dmem_n37, mem_stage_inst_dmem_n36,
         mem_stage_inst_dmem_n35, mem_stage_inst_dmem_n34,
         mem_stage_inst_dmem_n33, mem_stage_inst_dmem_n32,
         mem_stage_inst_dmem_n31, mem_stage_inst_dmem_n30,
         mem_stage_inst_dmem_n29, mem_stage_inst_dmem_n28,
         mem_stage_inst_dmem_n27, mem_stage_inst_dmem_n26,
         mem_stage_inst_dmem_n25, mem_stage_inst_dmem_n24,
         mem_stage_inst_dmem_n23, mem_stage_inst_dmem_n22,
         mem_stage_inst_dmem_n21, mem_stage_inst_dmem_n20,
         mem_stage_inst_dmem_n19, mem_stage_inst_dmem_n18,
         mem_stage_inst_dmem_n17, mem_stage_inst_dmem_n16,
         mem_stage_inst_dmem_n15, mem_stage_inst_dmem_n14,
         mem_stage_inst_dmem_n13, mem_stage_inst_dmem_n12,
         mem_stage_inst_dmem_n11, mem_stage_inst_dmem_n10,
         mem_stage_inst_dmem_n9, mem_stage_inst_dmem_n8,
         mem_stage_inst_dmem_n7, mem_stage_inst_dmem_n6,
         mem_stage_inst_dmem_n5, mem_stage_inst_dmem_n4,
         mem_stage_inst_dmem_n3, mem_stage_inst_dmem_n2,
         mem_stage_inst_dmem_n1, mem_stage_inst_dmem_n4660,
         mem_stage_inst_dmem_n4659, mem_stage_inst_dmem_n4658,
         mem_stage_inst_dmem_n4657, mem_stage_inst_dmem_n4656,
         mem_stage_inst_dmem_n4655, mem_stage_inst_dmem_n4654,
         mem_stage_inst_dmem_n4653, mem_stage_inst_dmem_n4652,
         mem_stage_inst_dmem_n4651, mem_stage_inst_dmem_n4650,
         mem_stage_inst_dmem_n4649, mem_stage_inst_dmem_n4648,
         mem_stage_inst_dmem_n4647, mem_stage_inst_dmem_n4646,
         mem_stage_inst_dmem_n4645, mem_stage_inst_dmem_n4644,
         mem_stage_inst_dmem_n4643, mem_stage_inst_dmem_n4642,
         mem_stage_inst_dmem_n4641, mem_stage_inst_dmem_n4640,
         mem_stage_inst_dmem_n4639, mem_stage_inst_dmem_n4638,
         mem_stage_inst_dmem_n4637, mem_stage_inst_dmem_n4636,
         mem_stage_inst_dmem_n4635, mem_stage_inst_dmem_n4634,
         mem_stage_inst_dmem_n4633, mem_stage_inst_dmem_n4632,
         mem_stage_inst_dmem_n4631, mem_stage_inst_dmem_n4630,
         mem_stage_inst_dmem_n4629, mem_stage_inst_dmem_n4628,
         mem_stage_inst_dmem_n4627, mem_stage_inst_dmem_n4626,
         mem_stage_inst_dmem_n4625, mem_stage_inst_dmem_n4624,
         mem_stage_inst_dmem_n4623, mem_stage_inst_dmem_n4622,
         mem_stage_inst_dmem_n4621, mem_stage_inst_dmem_n4620,
         mem_stage_inst_dmem_n4619, mem_stage_inst_dmem_n4618,
         mem_stage_inst_dmem_n4617, mem_stage_inst_dmem_n4616,
         mem_stage_inst_dmem_n4615, mem_stage_inst_dmem_n4614,
         mem_stage_inst_dmem_n4613, mem_stage_inst_dmem_n4612,
         mem_stage_inst_dmem_n4611, mem_stage_inst_dmem_n4610,
         mem_stage_inst_dmem_n4609, mem_stage_inst_dmem_n4608,
         mem_stage_inst_dmem_n4607, mem_stage_inst_dmem_n4606,
         mem_stage_inst_dmem_n4605, mem_stage_inst_dmem_n4604,
         mem_stage_inst_dmem_n4603, mem_stage_inst_dmem_n4602,
         mem_stage_inst_dmem_n4601, mem_stage_inst_dmem_n4600,
         mem_stage_inst_dmem_n4599, mem_stage_inst_dmem_n4598,
         mem_stage_inst_dmem_n4597, mem_stage_inst_dmem_n4596,
         mem_stage_inst_dmem_n4595, mem_stage_inst_dmem_n4594,
         mem_stage_inst_dmem_n4593, mem_stage_inst_dmem_n4592,
         mem_stage_inst_dmem_n4591, mem_stage_inst_dmem_n4590,
         mem_stage_inst_dmem_n4589, mem_stage_inst_dmem_n4588,
         mem_stage_inst_dmem_n4587, mem_stage_inst_dmem_n4586,
         mem_stage_inst_dmem_n4585, mem_stage_inst_dmem_n4584,
         mem_stage_inst_dmem_n4583, mem_stage_inst_dmem_n4582,
         mem_stage_inst_dmem_n4581, mem_stage_inst_dmem_n4580,
         mem_stage_inst_dmem_n4579, mem_stage_inst_dmem_n4578,
         mem_stage_inst_dmem_n4577, mem_stage_inst_dmem_n4576,
         mem_stage_inst_dmem_n4575, mem_stage_inst_dmem_n4574,
         mem_stage_inst_dmem_n4573, mem_stage_inst_dmem_n4572,
         mem_stage_inst_dmem_n4571, mem_stage_inst_dmem_n4570,
         mem_stage_inst_dmem_n4569, mem_stage_inst_dmem_n4568,
         mem_stage_inst_dmem_n4567, mem_stage_inst_dmem_n4566,
         mem_stage_inst_dmem_n4565, mem_stage_inst_dmem_n4564,
         mem_stage_inst_dmem_n4563, mem_stage_inst_dmem_n4562,
         mem_stage_inst_dmem_n4561, mem_stage_inst_dmem_n4560,
         mem_stage_inst_dmem_n4559, mem_stage_inst_dmem_n4558,
         mem_stage_inst_dmem_n4557, mem_stage_inst_dmem_n4556,
         mem_stage_inst_dmem_n4555, mem_stage_inst_dmem_n4554,
         mem_stage_inst_dmem_n4553, mem_stage_inst_dmem_n4552,
         mem_stage_inst_dmem_n4551, mem_stage_inst_dmem_n4550,
         mem_stage_inst_dmem_n4549, mem_stage_inst_dmem_n4548,
         mem_stage_inst_dmem_n4547, mem_stage_inst_dmem_n4546,
         mem_stage_inst_dmem_n4545, mem_stage_inst_dmem_n4544,
         mem_stage_inst_dmem_n4543, mem_stage_inst_dmem_n4542,
         mem_stage_inst_dmem_n4541, mem_stage_inst_dmem_n4540,
         mem_stage_inst_dmem_n4539, mem_stage_inst_dmem_n4538,
         mem_stage_inst_dmem_n4537, mem_stage_inst_dmem_n4536,
         mem_stage_inst_dmem_n4535, mem_stage_inst_dmem_n4534,
         mem_stage_inst_dmem_n4533, mem_stage_inst_dmem_n4532,
         mem_stage_inst_dmem_n4531, mem_stage_inst_dmem_n4530,
         mem_stage_inst_dmem_n4529, mem_stage_inst_dmem_n4528,
         mem_stage_inst_dmem_n4527, mem_stage_inst_dmem_n4526,
         mem_stage_inst_dmem_n4525, mem_stage_inst_dmem_n4524,
         mem_stage_inst_dmem_n4523, mem_stage_inst_dmem_n4522,
         mem_stage_inst_dmem_n4521, mem_stage_inst_dmem_n4520,
         mem_stage_inst_dmem_n4519, mem_stage_inst_dmem_n4518,
         mem_stage_inst_dmem_n4517, mem_stage_inst_dmem_n4516,
         mem_stage_inst_dmem_n4515, mem_stage_inst_dmem_n4514,
         mem_stage_inst_dmem_n4513, mem_stage_inst_dmem_n4512,
         mem_stage_inst_dmem_n4511, mem_stage_inst_dmem_n4510,
         mem_stage_inst_dmem_n4509, mem_stage_inst_dmem_n4508,
         mem_stage_inst_dmem_n4507, mem_stage_inst_dmem_n4506,
         mem_stage_inst_dmem_n4505, mem_stage_inst_dmem_n4504,
         mem_stage_inst_dmem_n4503, mem_stage_inst_dmem_n4502,
         mem_stage_inst_dmem_n4501, mem_stage_inst_dmem_n4500,
         mem_stage_inst_dmem_n4499, mem_stage_inst_dmem_n4498,
         mem_stage_inst_dmem_n4497, mem_stage_inst_dmem_n4496,
         mem_stage_inst_dmem_n4495, mem_stage_inst_dmem_n4494,
         mem_stage_inst_dmem_n4493, mem_stage_inst_dmem_n4492,
         mem_stage_inst_dmem_n4491, mem_stage_inst_dmem_n4490,
         mem_stage_inst_dmem_n4489, mem_stage_inst_dmem_n4488,
         mem_stage_inst_dmem_n4487, mem_stage_inst_dmem_n4486,
         mem_stage_inst_dmem_n4485, mem_stage_inst_dmem_n4484,
         mem_stage_inst_dmem_n4483, mem_stage_inst_dmem_n4482,
         mem_stage_inst_dmem_n4481, mem_stage_inst_dmem_n4480,
         mem_stage_inst_dmem_n4479, mem_stage_inst_dmem_n4478,
         mem_stage_inst_dmem_n4477, mem_stage_inst_dmem_n4476,
         mem_stage_inst_dmem_n4475, mem_stage_inst_dmem_n4474,
         mem_stage_inst_dmem_n4473, mem_stage_inst_dmem_n4472,
         mem_stage_inst_dmem_n4471, mem_stage_inst_dmem_n4470,
         mem_stage_inst_dmem_n4469, mem_stage_inst_dmem_n4468,
         mem_stage_inst_dmem_n4467, mem_stage_inst_dmem_n4466,
         mem_stage_inst_dmem_n4465, mem_stage_inst_dmem_n4464,
         mem_stage_inst_dmem_n4463, mem_stage_inst_dmem_n4462,
         mem_stage_inst_dmem_n4461, mem_stage_inst_dmem_n4460,
         mem_stage_inst_dmem_n4459, mem_stage_inst_dmem_n4458,
         mem_stage_inst_dmem_n4457, mem_stage_inst_dmem_n4456,
         mem_stage_inst_dmem_n4455, mem_stage_inst_dmem_n4454,
         mem_stage_inst_dmem_n4453, mem_stage_inst_dmem_n4452,
         mem_stage_inst_dmem_n4451, mem_stage_inst_dmem_n4450,
         mem_stage_inst_dmem_n4449, mem_stage_inst_dmem_n4448,
         mem_stage_inst_dmem_n4447, mem_stage_inst_dmem_n4446,
         mem_stage_inst_dmem_n4445, mem_stage_inst_dmem_n4444,
         mem_stage_inst_dmem_n4443, mem_stage_inst_dmem_n4442,
         mem_stage_inst_dmem_n4441, mem_stage_inst_dmem_n4440,
         mem_stage_inst_dmem_n4439, mem_stage_inst_dmem_n4438,
         mem_stage_inst_dmem_n4437, mem_stage_inst_dmem_n4436,
         mem_stage_inst_dmem_n4435, mem_stage_inst_dmem_n4434,
         mem_stage_inst_dmem_n4433, mem_stage_inst_dmem_n4432,
         mem_stage_inst_dmem_n4431, mem_stage_inst_dmem_n4430,
         mem_stage_inst_dmem_n4429, mem_stage_inst_dmem_n4428,
         mem_stage_inst_dmem_n4427, mem_stage_inst_dmem_n4426,
         mem_stage_inst_dmem_n4425, mem_stage_inst_dmem_n4424,
         mem_stage_inst_dmem_n4423, mem_stage_inst_dmem_n4422,
         mem_stage_inst_dmem_n4421, mem_stage_inst_dmem_n4420,
         mem_stage_inst_dmem_n4419, mem_stage_inst_dmem_n4418,
         mem_stage_inst_dmem_n4417, mem_stage_inst_dmem_n4416,
         mem_stage_inst_dmem_n4415, mem_stage_inst_dmem_n4414,
         mem_stage_inst_dmem_n4413, mem_stage_inst_dmem_n4412,
         mem_stage_inst_dmem_n4411, mem_stage_inst_dmem_n4410,
         mem_stage_inst_dmem_n4409, mem_stage_inst_dmem_n4408,
         mem_stage_inst_dmem_n4407, mem_stage_inst_dmem_n4406,
         mem_stage_inst_dmem_n4405, mem_stage_inst_dmem_n4404,
         mem_stage_inst_dmem_n4403, mem_stage_inst_dmem_n4402,
         mem_stage_inst_dmem_n4401, mem_stage_inst_dmem_n4400,
         mem_stage_inst_dmem_n4399, mem_stage_inst_dmem_n4398,
         mem_stage_inst_dmem_n4397, mem_stage_inst_dmem_n4396,
         mem_stage_inst_dmem_n4395, mem_stage_inst_dmem_n4394,
         mem_stage_inst_dmem_n4393, mem_stage_inst_dmem_n4392,
         mem_stage_inst_dmem_n4391, mem_stage_inst_dmem_n4390,
         mem_stage_inst_dmem_n4389, mem_stage_inst_dmem_n4388,
         mem_stage_inst_dmem_n4387, mem_stage_inst_dmem_n4386,
         mem_stage_inst_dmem_n4385, mem_stage_inst_dmem_n4384,
         mem_stage_inst_dmem_n4383, mem_stage_inst_dmem_n4382,
         mem_stage_inst_dmem_n4381, mem_stage_inst_dmem_n4380,
         mem_stage_inst_dmem_n4379, mem_stage_inst_dmem_n4378,
         mem_stage_inst_dmem_n4377, mem_stage_inst_dmem_n4376,
         mem_stage_inst_dmem_n4375, mem_stage_inst_dmem_n4374,
         mem_stage_inst_dmem_n4373, mem_stage_inst_dmem_n4372,
         mem_stage_inst_dmem_n4371, mem_stage_inst_dmem_n4370,
         mem_stage_inst_dmem_n4369, mem_stage_inst_dmem_n4368,
         mem_stage_inst_dmem_n4367, mem_stage_inst_dmem_n4366,
         mem_stage_inst_dmem_n4365, mem_stage_inst_dmem_n4364,
         mem_stage_inst_dmem_n4363, mem_stage_inst_dmem_n4362,
         mem_stage_inst_dmem_n4361, mem_stage_inst_dmem_n4360,
         mem_stage_inst_dmem_n4359, mem_stage_inst_dmem_n4358,
         mem_stage_inst_dmem_n4357, mem_stage_inst_dmem_n4356,
         mem_stage_inst_dmem_n4355, mem_stage_inst_dmem_n4354,
         mem_stage_inst_dmem_n4353, mem_stage_inst_dmem_n4352,
         mem_stage_inst_dmem_n4351, mem_stage_inst_dmem_n4350,
         mem_stage_inst_dmem_n4349, mem_stage_inst_dmem_n4348,
         mem_stage_inst_dmem_n4347, mem_stage_inst_dmem_n4346,
         mem_stage_inst_dmem_n4345, mem_stage_inst_dmem_n4344,
         mem_stage_inst_dmem_n4343, mem_stage_inst_dmem_n4342,
         mem_stage_inst_dmem_n4341, mem_stage_inst_dmem_n4340,
         mem_stage_inst_dmem_n4339, mem_stage_inst_dmem_n4338,
         mem_stage_inst_dmem_n4337, mem_stage_inst_dmem_n4336,
         mem_stage_inst_dmem_n4335, mem_stage_inst_dmem_n4334,
         mem_stage_inst_dmem_n4333, mem_stage_inst_dmem_n4332,
         mem_stage_inst_dmem_n4331, mem_stage_inst_dmem_n4330,
         mem_stage_inst_dmem_n4329, mem_stage_inst_dmem_n4328,
         mem_stage_inst_dmem_n4327, mem_stage_inst_dmem_n4326,
         mem_stage_inst_dmem_n4325, mem_stage_inst_dmem_n4324,
         mem_stage_inst_dmem_n4323, mem_stage_inst_dmem_n4322,
         mem_stage_inst_dmem_n4321, mem_stage_inst_dmem_n4320,
         mem_stage_inst_dmem_n4319, mem_stage_inst_dmem_n4318,
         mem_stage_inst_dmem_n4317, mem_stage_inst_dmem_n4316,
         mem_stage_inst_dmem_n4315, mem_stage_inst_dmem_n4314,
         mem_stage_inst_dmem_n4313, mem_stage_inst_dmem_n4312,
         mem_stage_inst_dmem_n4311, mem_stage_inst_dmem_n4310,
         mem_stage_inst_dmem_n4309, mem_stage_inst_dmem_n4308,
         mem_stage_inst_dmem_n4307, mem_stage_inst_dmem_n4306,
         mem_stage_inst_dmem_n4305, mem_stage_inst_dmem_n4304,
         mem_stage_inst_dmem_n4303, mem_stage_inst_dmem_n4302,
         mem_stage_inst_dmem_n4301, mem_stage_inst_dmem_n4300,
         mem_stage_inst_dmem_n4299, mem_stage_inst_dmem_n4298,
         mem_stage_inst_dmem_n4297, mem_stage_inst_dmem_n4296,
         mem_stage_inst_dmem_n4295, mem_stage_inst_dmem_n4294,
         mem_stage_inst_dmem_n4293, mem_stage_inst_dmem_n4292,
         mem_stage_inst_dmem_n4291, mem_stage_inst_dmem_n4290,
         mem_stage_inst_dmem_n4289, mem_stage_inst_dmem_n4288,
         mem_stage_inst_dmem_n4287, mem_stage_inst_dmem_n4286,
         mem_stage_inst_dmem_n4285, mem_stage_inst_dmem_n4284,
         mem_stage_inst_dmem_n4283, mem_stage_inst_dmem_n4282,
         mem_stage_inst_dmem_n4281, mem_stage_inst_dmem_n4280,
         mem_stage_inst_dmem_n4279, mem_stage_inst_dmem_n4278,
         mem_stage_inst_dmem_n4277, mem_stage_inst_dmem_n4276,
         mem_stage_inst_dmem_n4275, mem_stage_inst_dmem_n4274,
         mem_stage_inst_dmem_n4273, mem_stage_inst_dmem_n4272,
         mem_stage_inst_dmem_n4271, mem_stage_inst_dmem_n4270,
         mem_stage_inst_dmem_n4269, mem_stage_inst_dmem_n4268,
         mem_stage_inst_dmem_n4267, mem_stage_inst_dmem_n4266,
         mem_stage_inst_dmem_n4265, mem_stage_inst_dmem_n4264,
         mem_stage_inst_dmem_n4263, mem_stage_inst_dmem_n4262,
         mem_stage_inst_dmem_n4261, mem_stage_inst_dmem_n4260,
         mem_stage_inst_dmem_n4259, mem_stage_inst_dmem_n4258,
         mem_stage_inst_dmem_n4257, mem_stage_inst_dmem_n4256,
         mem_stage_inst_dmem_n4255, mem_stage_inst_dmem_n4254,
         mem_stage_inst_dmem_n4253, mem_stage_inst_dmem_n4252,
         mem_stage_inst_dmem_n4251, mem_stage_inst_dmem_n4250,
         mem_stage_inst_dmem_n4249, mem_stage_inst_dmem_n4248,
         mem_stage_inst_dmem_n4247, mem_stage_inst_dmem_n4246,
         mem_stage_inst_dmem_n4245, mem_stage_inst_dmem_n4244,
         mem_stage_inst_dmem_n4243, mem_stage_inst_dmem_n4242,
         mem_stage_inst_dmem_n4241, mem_stage_inst_dmem_n4240,
         mem_stage_inst_dmem_n4239, mem_stage_inst_dmem_n4238,
         mem_stage_inst_dmem_n4237, mem_stage_inst_dmem_n4236,
         mem_stage_inst_dmem_n4235, mem_stage_inst_dmem_n4234,
         mem_stage_inst_dmem_n4233, mem_stage_inst_dmem_n4232,
         mem_stage_inst_dmem_n4231, mem_stage_inst_dmem_n4230,
         mem_stage_inst_dmem_n4229, mem_stage_inst_dmem_n4228,
         mem_stage_inst_dmem_n4227, mem_stage_inst_dmem_n4226,
         mem_stage_inst_dmem_n4225, mem_stage_inst_dmem_n4224,
         mem_stage_inst_dmem_n4223, mem_stage_inst_dmem_n4222,
         mem_stage_inst_dmem_n4221, mem_stage_inst_dmem_n4220,
         mem_stage_inst_dmem_n4219, mem_stage_inst_dmem_n4218,
         mem_stage_inst_dmem_n4217, mem_stage_inst_dmem_n4216,
         mem_stage_inst_dmem_n4215, mem_stage_inst_dmem_n4214,
         mem_stage_inst_dmem_n4213, mem_stage_inst_dmem_n4212,
         mem_stage_inst_dmem_n4211, mem_stage_inst_dmem_n4210,
         mem_stage_inst_dmem_n4209, mem_stage_inst_dmem_n4208,
         mem_stage_inst_dmem_n4207, mem_stage_inst_dmem_n4206,
         mem_stage_inst_dmem_n4205, mem_stage_inst_dmem_n4204,
         mem_stage_inst_dmem_n4203, mem_stage_inst_dmem_n4202,
         mem_stage_inst_dmem_n4201, mem_stage_inst_dmem_n4200,
         mem_stage_inst_dmem_n4199, mem_stage_inst_dmem_n4198,
         mem_stage_inst_dmem_n4197, mem_stage_inst_dmem_n4196,
         mem_stage_inst_dmem_n4195, mem_stage_inst_dmem_n4194,
         mem_stage_inst_dmem_n4193, mem_stage_inst_dmem_n4192,
         mem_stage_inst_dmem_n4191, mem_stage_inst_dmem_n4190,
         mem_stage_inst_dmem_n4189, mem_stage_inst_dmem_n4188,
         mem_stage_inst_dmem_n4187, mem_stage_inst_dmem_n4186,
         mem_stage_inst_dmem_n4185, mem_stage_inst_dmem_n4184,
         mem_stage_inst_dmem_n4183, mem_stage_inst_dmem_n4182,
         mem_stage_inst_dmem_n4181, mem_stage_inst_dmem_n4180,
         mem_stage_inst_dmem_n4179, mem_stage_inst_dmem_n4178,
         mem_stage_inst_dmem_n4177, mem_stage_inst_dmem_n4176,
         mem_stage_inst_dmem_n4175, mem_stage_inst_dmem_n4174,
         mem_stage_inst_dmem_n4173, mem_stage_inst_dmem_n4172,
         mem_stage_inst_dmem_n4171, mem_stage_inst_dmem_n4170,
         mem_stage_inst_dmem_n4169, mem_stage_inst_dmem_n4168,
         mem_stage_inst_dmem_n4167, mem_stage_inst_dmem_n4166,
         mem_stage_inst_dmem_n4165, mem_stage_inst_dmem_n4164,
         mem_stage_inst_dmem_n4163, mem_stage_inst_dmem_n4162,
         mem_stage_inst_dmem_n4161, mem_stage_inst_dmem_n4160,
         mem_stage_inst_dmem_n4159, mem_stage_inst_dmem_n4158,
         mem_stage_inst_dmem_n4157, mem_stage_inst_dmem_n4156,
         mem_stage_inst_dmem_n4155, mem_stage_inst_dmem_n4154,
         mem_stage_inst_dmem_n4153, mem_stage_inst_dmem_n4152,
         mem_stage_inst_dmem_n4151, mem_stage_inst_dmem_n4150,
         mem_stage_inst_dmem_n4149, mem_stage_inst_dmem_n4148,
         mem_stage_inst_dmem_n4147, mem_stage_inst_dmem_n4146,
         mem_stage_inst_dmem_n4145, mem_stage_inst_dmem_n4144,
         mem_stage_inst_dmem_n4143, mem_stage_inst_dmem_n4142,
         mem_stage_inst_dmem_n4141, mem_stage_inst_dmem_n4140,
         mem_stage_inst_dmem_n4139, mem_stage_inst_dmem_n4138,
         mem_stage_inst_dmem_n4137, mem_stage_inst_dmem_n4136,
         mem_stage_inst_dmem_n4135, mem_stage_inst_dmem_n4134,
         mem_stage_inst_dmem_n4133, mem_stage_inst_dmem_n4132,
         mem_stage_inst_dmem_n4131, mem_stage_inst_dmem_n4130,
         mem_stage_inst_dmem_n4129, mem_stage_inst_dmem_n4128,
         mem_stage_inst_dmem_n4127, mem_stage_inst_dmem_n4126,
         mem_stage_inst_dmem_n4125, mem_stage_inst_dmem_n4124,
         mem_stage_inst_dmem_n4123, mem_stage_inst_dmem_n4122,
         mem_stage_inst_dmem_n4121, mem_stage_inst_dmem_n4120,
         mem_stage_inst_dmem_n4119, mem_stage_inst_dmem_n4118,
         mem_stage_inst_dmem_n4117, mem_stage_inst_dmem_n4116,
         mem_stage_inst_dmem_n4115, mem_stage_inst_dmem_n4114,
         mem_stage_inst_dmem_n4113, mem_stage_inst_dmem_n4112,
         mem_stage_inst_dmem_n4111, mem_stage_inst_dmem_n4110,
         mem_stage_inst_dmem_n4109, mem_stage_inst_dmem_n4108,
         mem_stage_inst_dmem_n4107, mem_stage_inst_dmem_n4106,
         mem_stage_inst_dmem_n4105, mem_stage_inst_dmem_n4104,
         mem_stage_inst_dmem_n4103, mem_stage_inst_dmem_n4102,
         mem_stage_inst_dmem_n4101, mem_stage_inst_dmem_n4100,
         mem_stage_inst_dmem_n4099, mem_stage_inst_dmem_n4098,
         mem_stage_inst_dmem_n4097, mem_stage_inst_dmem_n4096,
         mem_stage_inst_dmem_n4095, mem_stage_inst_dmem_n4094,
         mem_stage_inst_dmem_n4093, mem_stage_inst_dmem_n4092,
         mem_stage_inst_dmem_n4091, mem_stage_inst_dmem_n4090,
         mem_stage_inst_dmem_n4089, mem_stage_inst_dmem_n4088,
         mem_stage_inst_dmem_n4087, mem_stage_inst_dmem_n4086,
         mem_stage_inst_dmem_n4085, mem_stage_inst_dmem_n4084,
         mem_stage_inst_dmem_n4083, mem_stage_inst_dmem_n4082,
         mem_stage_inst_dmem_n4081, mem_stage_inst_dmem_n4080,
         mem_stage_inst_dmem_n4079, mem_stage_inst_dmem_n4078,
         mem_stage_inst_dmem_n4077, mem_stage_inst_dmem_n4076,
         mem_stage_inst_dmem_n4075, mem_stage_inst_dmem_n4074,
         mem_stage_inst_dmem_n4073, mem_stage_inst_dmem_n4072,
         mem_stage_inst_dmem_n4071, mem_stage_inst_dmem_n4070,
         mem_stage_inst_dmem_n4069, mem_stage_inst_dmem_n4068,
         mem_stage_inst_dmem_n4067, mem_stage_inst_dmem_n4066,
         mem_stage_inst_dmem_n4065, mem_stage_inst_dmem_n4064,
         mem_stage_inst_dmem_n4063, mem_stage_inst_dmem_n4062,
         mem_stage_inst_dmem_n4061, mem_stage_inst_dmem_n4060,
         mem_stage_inst_dmem_n4059, mem_stage_inst_dmem_n4058,
         mem_stage_inst_dmem_n4057, mem_stage_inst_dmem_n4056,
         mem_stage_inst_dmem_n4055, mem_stage_inst_dmem_n4054,
         mem_stage_inst_dmem_n4053, mem_stage_inst_dmem_n4052,
         mem_stage_inst_dmem_n4051, mem_stage_inst_dmem_n4050,
         mem_stage_inst_dmem_n4049, mem_stage_inst_dmem_n4048,
         mem_stage_inst_dmem_n4047, mem_stage_inst_dmem_n4046,
         mem_stage_inst_dmem_n4045, mem_stage_inst_dmem_n4044,
         mem_stage_inst_dmem_n4043, mem_stage_inst_dmem_n4042,
         mem_stage_inst_dmem_n4041, mem_stage_inst_dmem_n4040,
         mem_stage_inst_dmem_n4039, mem_stage_inst_dmem_n4038,
         mem_stage_inst_dmem_n4037, mem_stage_inst_dmem_n4036,
         mem_stage_inst_dmem_n4035, mem_stage_inst_dmem_n4034,
         mem_stage_inst_dmem_n4033, mem_stage_inst_dmem_n4032,
         mem_stage_inst_dmem_n4031, mem_stage_inst_dmem_n4030,
         mem_stage_inst_dmem_n4029, mem_stage_inst_dmem_n4028,
         mem_stage_inst_dmem_n4027, mem_stage_inst_dmem_n4026,
         mem_stage_inst_dmem_n4025, mem_stage_inst_dmem_n4024,
         mem_stage_inst_dmem_n4023, mem_stage_inst_dmem_n4022,
         mem_stage_inst_dmem_n4021, mem_stage_inst_dmem_n4020,
         mem_stage_inst_dmem_n4019, mem_stage_inst_dmem_n4018,
         mem_stage_inst_dmem_n4017, mem_stage_inst_dmem_n4016,
         mem_stage_inst_dmem_n4015, mem_stage_inst_dmem_n4014,
         mem_stage_inst_dmem_n4013, mem_stage_inst_dmem_n4012,
         mem_stage_inst_dmem_n4011, mem_stage_inst_dmem_n4010,
         mem_stage_inst_dmem_n4009, mem_stage_inst_dmem_n4008,
         mem_stage_inst_dmem_n4007, mem_stage_inst_dmem_n4006,
         mem_stage_inst_dmem_n4005, mem_stage_inst_dmem_n4004,
         mem_stage_inst_dmem_n4003, mem_stage_inst_dmem_n4002,
         mem_stage_inst_dmem_n4001, mem_stage_inst_dmem_n4000,
         mem_stage_inst_dmem_n3999, mem_stage_inst_dmem_n3998,
         mem_stage_inst_dmem_n3997, mem_stage_inst_dmem_n3996,
         mem_stage_inst_dmem_n3995, mem_stage_inst_dmem_n3994,
         mem_stage_inst_dmem_n3993, mem_stage_inst_dmem_n3992,
         mem_stage_inst_dmem_n3991, mem_stage_inst_dmem_n3990,
         mem_stage_inst_dmem_n3989, mem_stage_inst_dmem_n3988,
         mem_stage_inst_dmem_n3987, mem_stage_inst_dmem_n3986,
         mem_stage_inst_dmem_n3985, mem_stage_inst_dmem_n3984,
         mem_stage_inst_dmem_n3983, mem_stage_inst_dmem_n3982,
         mem_stage_inst_dmem_n3981, mem_stage_inst_dmem_n3980,
         mem_stage_inst_dmem_n3979, mem_stage_inst_dmem_n3978,
         mem_stage_inst_dmem_n3977, mem_stage_inst_dmem_n3976,
         mem_stage_inst_dmem_n3975, mem_stage_inst_dmem_n3974,
         mem_stage_inst_dmem_n3973, mem_stage_inst_dmem_n3972,
         mem_stage_inst_dmem_n3971, mem_stage_inst_dmem_n3970,
         mem_stage_inst_dmem_n3969, mem_stage_inst_dmem_n3968,
         mem_stage_inst_dmem_n3967, mem_stage_inst_dmem_n3966,
         mem_stage_inst_dmem_n3965, mem_stage_inst_dmem_n3964,
         mem_stage_inst_dmem_n3963, mem_stage_inst_dmem_n3962,
         mem_stage_inst_dmem_n3961, mem_stage_inst_dmem_n3960,
         mem_stage_inst_dmem_n3959, mem_stage_inst_dmem_n3958,
         mem_stage_inst_dmem_n3957, mem_stage_inst_dmem_n3956,
         mem_stage_inst_dmem_n3955, mem_stage_inst_dmem_n3954,
         mem_stage_inst_dmem_n3953, mem_stage_inst_dmem_n3952,
         mem_stage_inst_dmem_n3951, mem_stage_inst_dmem_n3950,
         mem_stage_inst_dmem_n3949, mem_stage_inst_dmem_n3948,
         mem_stage_inst_dmem_n3947, mem_stage_inst_dmem_n3946,
         mem_stage_inst_dmem_n3945, mem_stage_inst_dmem_n3944,
         mem_stage_inst_dmem_n3943, mem_stage_inst_dmem_n3942,
         mem_stage_inst_dmem_n3941, mem_stage_inst_dmem_n3940,
         mem_stage_inst_dmem_n3939, mem_stage_inst_dmem_n3938,
         mem_stage_inst_dmem_n3937, mem_stage_inst_dmem_n3936,
         mem_stage_inst_dmem_n3935, mem_stage_inst_dmem_n3934,
         mem_stage_inst_dmem_n3933, mem_stage_inst_dmem_n3932,
         mem_stage_inst_dmem_n3931, mem_stage_inst_dmem_n3930,
         mem_stage_inst_dmem_n3929, mem_stage_inst_dmem_n3928,
         mem_stage_inst_dmem_n3927, mem_stage_inst_dmem_n3926,
         mem_stage_inst_dmem_n3925, mem_stage_inst_dmem_n3924,
         mem_stage_inst_dmem_n3923, mem_stage_inst_dmem_n3922,
         mem_stage_inst_dmem_n3921, mem_stage_inst_dmem_n3920,
         mem_stage_inst_dmem_n3919, mem_stage_inst_dmem_n3918,
         mem_stage_inst_dmem_n3917, mem_stage_inst_dmem_n3916,
         mem_stage_inst_dmem_n3915, mem_stage_inst_dmem_n3914,
         mem_stage_inst_dmem_n3913, mem_stage_inst_dmem_n3912,
         mem_stage_inst_dmem_n3911, mem_stage_inst_dmem_n3910,
         mem_stage_inst_dmem_n3909, mem_stage_inst_dmem_n3908,
         mem_stage_inst_dmem_n3907, mem_stage_inst_dmem_n3906,
         mem_stage_inst_dmem_n3905, mem_stage_inst_dmem_n3904,
         mem_stage_inst_dmem_n3903, mem_stage_inst_dmem_n3902,
         mem_stage_inst_dmem_n3901, mem_stage_inst_dmem_n3900,
         mem_stage_inst_dmem_n3899, mem_stage_inst_dmem_n3898,
         mem_stage_inst_dmem_n3897, mem_stage_inst_dmem_n3896,
         mem_stage_inst_dmem_n3895, mem_stage_inst_dmem_n3894,
         mem_stage_inst_dmem_n3893, mem_stage_inst_dmem_n3892,
         mem_stage_inst_dmem_n3891, mem_stage_inst_dmem_n3890,
         mem_stage_inst_dmem_n3889, mem_stage_inst_dmem_n3888,
         mem_stage_inst_dmem_n3887, mem_stage_inst_dmem_n3886,
         mem_stage_inst_dmem_n3885, mem_stage_inst_dmem_n3884,
         mem_stage_inst_dmem_n3883, mem_stage_inst_dmem_n3882,
         mem_stage_inst_dmem_n3881, mem_stage_inst_dmem_n3880,
         mem_stage_inst_dmem_n3879, mem_stage_inst_dmem_n3878,
         mem_stage_inst_dmem_n3877, mem_stage_inst_dmem_n3876,
         mem_stage_inst_dmem_n3875, mem_stage_inst_dmem_n3874,
         mem_stage_inst_dmem_n3873, mem_stage_inst_dmem_n3872,
         mem_stage_inst_dmem_n3871, mem_stage_inst_dmem_n3870,
         mem_stage_inst_dmem_n3869, mem_stage_inst_dmem_n3868,
         mem_stage_inst_dmem_n3867, mem_stage_inst_dmem_n3866,
         mem_stage_inst_dmem_n3865, mem_stage_inst_dmem_n3864,
         mem_stage_inst_dmem_n3863, mem_stage_inst_dmem_n3862,
         mem_stage_inst_dmem_n3861, mem_stage_inst_dmem_n3860,
         mem_stage_inst_dmem_n3859, mem_stage_inst_dmem_n3858,
         mem_stage_inst_dmem_n3857, mem_stage_inst_dmem_n3856,
         mem_stage_inst_dmem_n3855, mem_stage_inst_dmem_n3854,
         mem_stage_inst_dmem_n3853, mem_stage_inst_dmem_n3852,
         mem_stage_inst_dmem_n3851, mem_stage_inst_dmem_n3850,
         mem_stage_inst_dmem_n3849, mem_stage_inst_dmem_n3848,
         mem_stage_inst_dmem_n3847, mem_stage_inst_dmem_n3846,
         mem_stage_inst_dmem_n3845, mem_stage_inst_dmem_n3844,
         mem_stage_inst_dmem_n3843, mem_stage_inst_dmem_n3842,
         mem_stage_inst_dmem_n3841, mem_stage_inst_dmem_n3840,
         mem_stage_inst_dmem_n3839, mem_stage_inst_dmem_n3838,
         mem_stage_inst_dmem_n3837, mem_stage_inst_dmem_n3836,
         mem_stage_inst_dmem_n3835, mem_stage_inst_dmem_n3834,
         mem_stage_inst_dmem_n3833, mem_stage_inst_dmem_n3832,
         mem_stage_inst_dmem_n3831, mem_stage_inst_dmem_n3830,
         mem_stage_inst_dmem_n3829, mem_stage_inst_dmem_n3828,
         mem_stage_inst_dmem_n3827, mem_stage_inst_dmem_n3826,
         mem_stage_inst_dmem_n3825, mem_stage_inst_dmem_n3824,
         mem_stage_inst_dmem_n3823, mem_stage_inst_dmem_n3822,
         mem_stage_inst_dmem_n3821, mem_stage_inst_dmem_n3820,
         mem_stage_inst_dmem_n3819, mem_stage_inst_dmem_n3818,
         mem_stage_inst_dmem_n3817, mem_stage_inst_dmem_n3816,
         mem_stage_inst_dmem_n3815, mem_stage_inst_dmem_n3814,
         mem_stage_inst_dmem_n3813, mem_stage_inst_dmem_n3812,
         mem_stage_inst_dmem_n3811, mem_stage_inst_dmem_n3810,
         mem_stage_inst_dmem_n3809, mem_stage_inst_dmem_n3808,
         mem_stage_inst_dmem_n3807, mem_stage_inst_dmem_n3806,
         mem_stage_inst_dmem_n3805, mem_stage_inst_dmem_n3804,
         mem_stage_inst_dmem_n3803, mem_stage_inst_dmem_n3802,
         mem_stage_inst_dmem_n3801, mem_stage_inst_dmem_n3800,
         mem_stage_inst_dmem_n3799, mem_stage_inst_dmem_n3798,
         mem_stage_inst_dmem_n3797, mem_stage_inst_dmem_n3796,
         mem_stage_inst_dmem_n3795, mem_stage_inst_dmem_n3794,
         mem_stage_inst_dmem_n3793, mem_stage_inst_dmem_n3792,
         mem_stage_inst_dmem_n3791, mem_stage_inst_dmem_n3790,
         mem_stage_inst_dmem_n3789, mem_stage_inst_dmem_n3788,
         mem_stage_inst_dmem_n3787, mem_stage_inst_dmem_n3786,
         mem_stage_inst_dmem_n3785, mem_stage_inst_dmem_n3784,
         mem_stage_inst_dmem_n3783, mem_stage_inst_dmem_n3782,
         mem_stage_inst_dmem_n3781, mem_stage_inst_dmem_n3780,
         mem_stage_inst_dmem_n3779, mem_stage_inst_dmem_n3778,
         mem_stage_inst_dmem_n3777, mem_stage_inst_dmem_n3776,
         mem_stage_inst_dmem_n3775, mem_stage_inst_dmem_n3774,
         mem_stage_inst_dmem_n3773, mem_stage_inst_dmem_n3772,
         mem_stage_inst_dmem_n3771, mem_stage_inst_dmem_n3770,
         mem_stage_inst_dmem_n3769, mem_stage_inst_dmem_n3768,
         mem_stage_inst_dmem_n3767, mem_stage_inst_dmem_n3766,
         mem_stage_inst_dmem_n3765, mem_stage_inst_dmem_n3764,
         mem_stage_inst_dmem_n3763, mem_stage_inst_dmem_n3762,
         mem_stage_inst_dmem_n3761, mem_stage_inst_dmem_n3760,
         mem_stage_inst_dmem_n3759, mem_stage_inst_dmem_n3758,
         mem_stage_inst_dmem_n3757, mem_stage_inst_dmem_n3756,
         mem_stage_inst_dmem_n3755, mem_stage_inst_dmem_n3754,
         mem_stage_inst_dmem_n3753, mem_stage_inst_dmem_n3752,
         mem_stage_inst_dmem_n3751, mem_stage_inst_dmem_n3750,
         mem_stage_inst_dmem_n3749, mem_stage_inst_dmem_n3748,
         mem_stage_inst_dmem_n3747, mem_stage_inst_dmem_n3746,
         mem_stage_inst_dmem_n3745, mem_stage_inst_dmem_n3744,
         mem_stage_inst_dmem_n3743, mem_stage_inst_dmem_n3742,
         mem_stage_inst_dmem_n3741, mem_stage_inst_dmem_n3740,
         mem_stage_inst_dmem_n3739, mem_stage_inst_dmem_n3738,
         mem_stage_inst_dmem_n3737, mem_stage_inst_dmem_n3736,
         mem_stage_inst_dmem_n3735, mem_stage_inst_dmem_n3734,
         mem_stage_inst_dmem_n3733, mem_stage_inst_dmem_n3732,
         mem_stage_inst_dmem_n3731, mem_stage_inst_dmem_n3730,
         mem_stage_inst_dmem_n3729, mem_stage_inst_dmem_n3728,
         mem_stage_inst_dmem_n3727, mem_stage_inst_dmem_n3726,
         mem_stage_inst_dmem_n3725, mem_stage_inst_dmem_n3724,
         mem_stage_inst_dmem_n3723, mem_stage_inst_dmem_n3722,
         mem_stage_inst_dmem_n3721, mem_stage_inst_dmem_n3720,
         mem_stage_inst_dmem_n3719, mem_stage_inst_dmem_n3718,
         mem_stage_inst_dmem_n3717, mem_stage_inst_dmem_n3716,
         mem_stage_inst_dmem_n3715, mem_stage_inst_dmem_n3714,
         mem_stage_inst_dmem_n3713, mem_stage_inst_dmem_n3712,
         mem_stage_inst_dmem_n3711, mem_stage_inst_dmem_n3710,
         mem_stage_inst_dmem_n3709, mem_stage_inst_dmem_n3708,
         mem_stage_inst_dmem_n3707, mem_stage_inst_dmem_n3706,
         mem_stage_inst_dmem_n3705, mem_stage_inst_dmem_n3704,
         mem_stage_inst_dmem_n3703, mem_stage_inst_dmem_n3702,
         mem_stage_inst_dmem_n3701, mem_stage_inst_dmem_n3700,
         mem_stage_inst_dmem_n3699, mem_stage_inst_dmem_n3698,
         mem_stage_inst_dmem_n3697, mem_stage_inst_dmem_n3696,
         mem_stage_inst_dmem_n3695, mem_stage_inst_dmem_n3694,
         mem_stage_inst_dmem_n3693, mem_stage_inst_dmem_n3692,
         mem_stage_inst_dmem_n3691, mem_stage_inst_dmem_n3690,
         mem_stage_inst_dmem_n3689, mem_stage_inst_dmem_n3688,
         mem_stage_inst_dmem_n3687, mem_stage_inst_dmem_n3686,
         mem_stage_inst_dmem_n3685, mem_stage_inst_dmem_n3684,
         mem_stage_inst_dmem_n3683, mem_stage_inst_dmem_n3682,
         mem_stage_inst_dmem_n3681, mem_stage_inst_dmem_n3680,
         mem_stage_inst_dmem_n3679, mem_stage_inst_dmem_n3678,
         mem_stage_inst_dmem_n3677, mem_stage_inst_dmem_n3676,
         mem_stage_inst_dmem_n3675, mem_stage_inst_dmem_n3674,
         mem_stage_inst_dmem_n3673, mem_stage_inst_dmem_n3672,
         mem_stage_inst_dmem_n3671, mem_stage_inst_dmem_n3670,
         mem_stage_inst_dmem_n3669, mem_stage_inst_dmem_n3668,
         mem_stage_inst_dmem_n3667, mem_stage_inst_dmem_n3666,
         mem_stage_inst_dmem_n3665, mem_stage_inst_dmem_n3664,
         mem_stage_inst_dmem_n3663, mem_stage_inst_dmem_n3662,
         mem_stage_inst_dmem_n3661, mem_stage_inst_dmem_n3660,
         mem_stage_inst_dmem_n3659, mem_stage_inst_dmem_n3658,
         mem_stage_inst_dmem_n3657, mem_stage_inst_dmem_n3656,
         mem_stage_inst_dmem_n3655, mem_stage_inst_dmem_n3654,
         mem_stage_inst_dmem_n3653, mem_stage_inst_dmem_n3652,
         mem_stage_inst_dmem_n3651, mem_stage_inst_dmem_n3650,
         mem_stage_inst_dmem_n3649, mem_stage_inst_dmem_n3648,
         mem_stage_inst_dmem_n3647, mem_stage_inst_dmem_n3646,
         mem_stage_inst_dmem_n3645, mem_stage_inst_dmem_n3644,
         mem_stage_inst_dmem_n3643, mem_stage_inst_dmem_n3642,
         mem_stage_inst_dmem_n3641, mem_stage_inst_dmem_n3640,
         mem_stage_inst_dmem_n3639, mem_stage_inst_dmem_n3638,
         mem_stage_inst_dmem_n3637, mem_stage_inst_dmem_n3636,
         mem_stage_inst_dmem_n3635, mem_stage_inst_dmem_n3634,
         mem_stage_inst_dmem_n3633, mem_stage_inst_dmem_n3632,
         mem_stage_inst_dmem_n3631, mem_stage_inst_dmem_n3630,
         mem_stage_inst_dmem_n3629, mem_stage_inst_dmem_n3628,
         mem_stage_inst_dmem_n3627, mem_stage_inst_dmem_n3626,
         mem_stage_inst_dmem_n3625, mem_stage_inst_dmem_n3624,
         mem_stage_inst_dmem_n3623, mem_stage_inst_dmem_n3622,
         mem_stage_inst_dmem_n3621, mem_stage_inst_dmem_n3620,
         mem_stage_inst_dmem_n3619, mem_stage_inst_dmem_n3618,
         mem_stage_inst_dmem_n3617, mem_stage_inst_dmem_n3616,
         mem_stage_inst_dmem_n3615, mem_stage_inst_dmem_n3614,
         mem_stage_inst_dmem_n3613, mem_stage_inst_dmem_n3612,
         mem_stage_inst_dmem_n3611, mem_stage_inst_dmem_n3610,
         mem_stage_inst_dmem_n3609, mem_stage_inst_dmem_n3608,
         mem_stage_inst_dmem_n3607, mem_stage_inst_dmem_n3606,
         mem_stage_inst_dmem_n3605, mem_stage_inst_dmem_n3604,
         mem_stage_inst_dmem_n3603, mem_stage_inst_dmem_n3602,
         mem_stage_inst_dmem_n3601, mem_stage_inst_dmem_n3600,
         mem_stage_inst_dmem_n3599, mem_stage_inst_dmem_n3598,
         mem_stage_inst_dmem_n3597, mem_stage_inst_dmem_n3596,
         mem_stage_inst_dmem_n3595, mem_stage_inst_dmem_n3594,
         mem_stage_inst_dmem_n3593, mem_stage_inst_dmem_n3592,
         mem_stage_inst_dmem_n3591, mem_stage_inst_dmem_n3590,
         mem_stage_inst_dmem_n3589, mem_stage_inst_dmem_n3588,
         mem_stage_inst_dmem_n3587, mem_stage_inst_dmem_n3586,
         mem_stage_inst_dmem_n3585, mem_stage_inst_dmem_n3584,
         mem_stage_inst_dmem_n3583, mem_stage_inst_dmem_n3582,
         mem_stage_inst_dmem_n3581, mem_stage_inst_dmem_n3580,
         mem_stage_inst_dmem_n3579, mem_stage_inst_dmem_n3578,
         mem_stage_inst_dmem_n3577, mem_stage_inst_dmem_n3576,
         mem_stage_inst_dmem_n3575, mem_stage_inst_dmem_n3574,
         mem_stage_inst_dmem_n3573, mem_stage_inst_dmem_n3572,
         mem_stage_inst_dmem_n3571, mem_stage_inst_dmem_n3570,
         mem_stage_inst_dmem_n3569, mem_stage_inst_dmem_n3568,
         mem_stage_inst_dmem_n3567, mem_stage_inst_dmem_n3566,
         mem_stage_inst_dmem_n3565, mem_stage_inst_dmem_n3564,
         mem_stage_inst_dmem_n3563, mem_stage_inst_dmem_n3562,
         mem_stage_inst_dmem_n3561, mem_stage_inst_dmem_n3560,
         mem_stage_inst_dmem_n3559, mem_stage_inst_dmem_n3558,
         mem_stage_inst_dmem_n3557, mem_stage_inst_dmem_n3556,
         mem_stage_inst_dmem_n3555, mem_stage_inst_dmem_n3554,
         mem_stage_inst_dmem_n3553, mem_stage_inst_dmem_n3552,
         mem_stage_inst_dmem_n3551, mem_stage_inst_dmem_n3550,
         mem_stage_inst_dmem_n3549, mem_stage_inst_dmem_n3548,
         mem_stage_inst_dmem_n3547, mem_stage_inst_dmem_n3546,
         mem_stage_inst_dmem_n3545, mem_stage_inst_dmem_n3544,
         mem_stage_inst_dmem_n3543, mem_stage_inst_dmem_n3542,
         mem_stage_inst_dmem_n3541, mem_stage_inst_dmem_n3540,
         mem_stage_inst_dmem_n3539, mem_stage_inst_dmem_n3538,
         mem_stage_inst_dmem_n3537, mem_stage_inst_dmem_n3536,
         mem_stage_inst_dmem_n3535, mem_stage_inst_dmem_n3534,
         mem_stage_inst_dmem_n3533, mem_stage_inst_dmem_n3532,
         mem_stage_inst_dmem_n3531, mem_stage_inst_dmem_n3530,
         mem_stage_inst_dmem_n3529, mem_stage_inst_dmem_n3528,
         mem_stage_inst_dmem_n3527, mem_stage_inst_dmem_n3526,
         mem_stage_inst_dmem_n3525, mem_stage_inst_dmem_n3524,
         mem_stage_inst_dmem_n3523, mem_stage_inst_dmem_n3522,
         mem_stage_inst_dmem_n3521, mem_stage_inst_dmem_n3520,
         mem_stage_inst_dmem_n3519, mem_stage_inst_dmem_n3518,
         mem_stage_inst_dmem_n3517, mem_stage_inst_dmem_n3516,
         mem_stage_inst_dmem_n3515, mem_stage_inst_dmem_n3514,
         mem_stage_inst_dmem_n3513, mem_stage_inst_dmem_n3512,
         mem_stage_inst_dmem_n3511, mem_stage_inst_dmem_n3510,
         mem_stage_inst_dmem_n3509, mem_stage_inst_dmem_n3508,
         mem_stage_inst_dmem_n3507, mem_stage_inst_dmem_n3506,
         mem_stage_inst_dmem_n3505, mem_stage_inst_dmem_n3504,
         mem_stage_inst_dmem_n3503, mem_stage_inst_dmem_n3502,
         mem_stage_inst_dmem_n3501, mem_stage_inst_dmem_n3500,
         mem_stage_inst_dmem_n3499, mem_stage_inst_dmem_n3498,
         mem_stage_inst_dmem_n3497, mem_stage_inst_dmem_n3496,
         mem_stage_inst_dmem_n3495, mem_stage_inst_dmem_n3494,
         mem_stage_inst_dmem_n3493, mem_stage_inst_dmem_n3492,
         mem_stage_inst_dmem_n3491, mem_stage_inst_dmem_n3490,
         mem_stage_inst_dmem_n3489, mem_stage_inst_dmem_n3488,
         mem_stage_inst_dmem_n3487, mem_stage_inst_dmem_n3486,
         mem_stage_inst_dmem_n3485, mem_stage_inst_dmem_n3484,
         mem_stage_inst_dmem_n3483, mem_stage_inst_dmem_n3482,
         mem_stage_inst_dmem_n3481, mem_stage_inst_dmem_n3480,
         mem_stage_inst_dmem_n3479, mem_stage_inst_dmem_n3478,
         mem_stage_inst_dmem_n3477, mem_stage_inst_dmem_n3476,
         mem_stage_inst_dmem_n3475, mem_stage_inst_dmem_n3474,
         mem_stage_inst_dmem_n3473, mem_stage_inst_dmem_n3472,
         mem_stage_inst_dmem_n3471, mem_stage_inst_dmem_n3470,
         mem_stage_inst_dmem_n3469, mem_stage_inst_dmem_n3468,
         mem_stage_inst_dmem_n3467, mem_stage_inst_dmem_n3466,
         mem_stage_inst_dmem_n3465, mem_stage_inst_dmem_n3464,
         mem_stage_inst_dmem_n3463, mem_stage_inst_dmem_n3462,
         mem_stage_inst_dmem_n3461, mem_stage_inst_dmem_n3460,
         mem_stage_inst_dmem_n3459, mem_stage_inst_dmem_n3458,
         mem_stage_inst_dmem_n3457, mem_stage_inst_dmem_n3456,
         mem_stage_inst_dmem_n3455, mem_stage_inst_dmem_n3454,
         mem_stage_inst_dmem_n3453, mem_stage_inst_dmem_n3452,
         mem_stage_inst_dmem_n3451, mem_stage_inst_dmem_n3450,
         mem_stage_inst_dmem_n3449, mem_stage_inst_dmem_n3448,
         mem_stage_inst_dmem_n3447, mem_stage_inst_dmem_n3446,
         mem_stage_inst_dmem_n3445, mem_stage_inst_dmem_n3444,
         mem_stage_inst_dmem_n3443, mem_stage_inst_dmem_n3442,
         mem_stage_inst_dmem_n3441, mem_stage_inst_dmem_n3440,
         mem_stage_inst_dmem_n3439, mem_stage_inst_dmem_n3438,
         mem_stage_inst_dmem_n3437, mem_stage_inst_dmem_n3436,
         mem_stage_inst_dmem_n3435, mem_stage_inst_dmem_n3434,
         mem_stage_inst_dmem_n3433, mem_stage_inst_dmem_n3432,
         mem_stage_inst_dmem_n3431, mem_stage_inst_dmem_n3430,
         mem_stage_inst_dmem_n3429, mem_stage_inst_dmem_n3428,
         mem_stage_inst_dmem_n3427, mem_stage_inst_dmem_n3426,
         mem_stage_inst_dmem_n3425, mem_stage_inst_dmem_n3424,
         mem_stage_inst_dmem_n3423, mem_stage_inst_dmem_n3422,
         mem_stage_inst_dmem_n3421, mem_stage_inst_dmem_n3420,
         mem_stage_inst_dmem_n3419, mem_stage_inst_dmem_n3418,
         mem_stage_inst_dmem_n3417, mem_stage_inst_dmem_n3416,
         mem_stage_inst_dmem_n3415, mem_stage_inst_dmem_n3414,
         mem_stage_inst_dmem_n3413, mem_stage_inst_dmem_n3412,
         mem_stage_inst_dmem_n3411, mem_stage_inst_dmem_n3410,
         mem_stage_inst_dmem_n3409, mem_stage_inst_dmem_n3408,
         mem_stage_inst_dmem_n3407, mem_stage_inst_dmem_n3406,
         mem_stage_inst_dmem_n3405, mem_stage_inst_dmem_n3404,
         mem_stage_inst_dmem_n3403, mem_stage_inst_dmem_n3402,
         mem_stage_inst_dmem_n3401, mem_stage_inst_dmem_n3400,
         mem_stage_inst_dmem_n3399, mem_stage_inst_dmem_n3398,
         mem_stage_inst_dmem_n3397, mem_stage_inst_dmem_n3396,
         mem_stage_inst_dmem_n3395, mem_stage_inst_dmem_n3394,
         mem_stage_inst_dmem_n3393, mem_stage_inst_dmem_n3392,
         mem_stage_inst_dmem_n3391, mem_stage_inst_dmem_n3390,
         mem_stage_inst_dmem_n3389, mem_stage_inst_dmem_n3388,
         mem_stage_inst_dmem_n3387, mem_stage_inst_dmem_n3386,
         mem_stage_inst_dmem_n3385, mem_stage_inst_dmem_n3384,
         mem_stage_inst_dmem_n3383, mem_stage_inst_dmem_n3382,
         mem_stage_inst_dmem_n3381, mem_stage_inst_dmem_n3380,
         mem_stage_inst_dmem_n3379, mem_stage_inst_dmem_n3378,
         mem_stage_inst_dmem_n3377, mem_stage_inst_dmem_n3376,
         mem_stage_inst_dmem_n3375, mem_stage_inst_dmem_n3374,
         mem_stage_inst_dmem_n3373, mem_stage_inst_dmem_n3372,
         mem_stage_inst_dmem_n3371, mem_stage_inst_dmem_n3370,
         mem_stage_inst_dmem_n3369, mem_stage_inst_dmem_n3368,
         mem_stage_inst_dmem_n3367, mem_stage_inst_dmem_n3366,
         mem_stage_inst_dmem_n3365, mem_stage_inst_dmem_n3364,
         mem_stage_inst_dmem_n3363, mem_stage_inst_dmem_n3362,
         mem_stage_inst_dmem_n3361, mem_stage_inst_dmem_n3360,
         mem_stage_inst_dmem_n3359, mem_stage_inst_dmem_n3358,
         mem_stage_inst_dmem_n3357, mem_stage_inst_dmem_n3356,
         mem_stage_inst_dmem_n3355, mem_stage_inst_dmem_n3354,
         mem_stage_inst_dmem_n3353, mem_stage_inst_dmem_n3352,
         mem_stage_inst_dmem_n3351, mem_stage_inst_dmem_n3350,
         mem_stage_inst_dmem_n3349, mem_stage_inst_dmem_n3348,
         mem_stage_inst_dmem_n3347, mem_stage_inst_dmem_n3346,
         mem_stage_inst_dmem_n3345, mem_stage_inst_dmem_n3344,
         mem_stage_inst_dmem_n3343, mem_stage_inst_dmem_n3342,
         mem_stage_inst_dmem_n3341, mem_stage_inst_dmem_n3340,
         mem_stage_inst_dmem_n3339, mem_stage_inst_dmem_n3338,
         mem_stage_inst_dmem_n3337, mem_stage_inst_dmem_n3336,
         mem_stage_inst_dmem_n3335, mem_stage_inst_dmem_n3334,
         mem_stage_inst_dmem_n3333, mem_stage_inst_dmem_n3332,
         mem_stage_inst_dmem_n3331, mem_stage_inst_dmem_n3330,
         mem_stage_inst_dmem_n3329, mem_stage_inst_dmem_n3328,
         mem_stage_inst_dmem_n3327, mem_stage_inst_dmem_n3326,
         mem_stage_inst_dmem_n3325, mem_stage_inst_dmem_n3324,
         mem_stage_inst_dmem_n3323, mem_stage_inst_dmem_n3322,
         mem_stage_inst_dmem_n3321, mem_stage_inst_dmem_n3320,
         mem_stage_inst_dmem_n3319, mem_stage_inst_dmem_n3318,
         mem_stage_inst_dmem_n3317, mem_stage_inst_dmem_n3316,
         mem_stage_inst_dmem_n3315, mem_stage_inst_dmem_n3314,
         mem_stage_inst_dmem_n3313, mem_stage_inst_dmem_n3312,
         mem_stage_inst_dmem_n3311, mem_stage_inst_dmem_n3310,
         mem_stage_inst_dmem_n3309, mem_stage_inst_dmem_n3308,
         mem_stage_inst_dmem_n3307, mem_stage_inst_dmem_n3306,
         mem_stage_inst_dmem_n3305, mem_stage_inst_dmem_n3304,
         mem_stage_inst_dmem_n3303, mem_stage_inst_dmem_n3302,
         mem_stage_inst_dmem_n3301, mem_stage_inst_dmem_n3300,
         mem_stage_inst_dmem_n3299, mem_stage_inst_dmem_n3298,
         mem_stage_inst_dmem_n3297, mem_stage_inst_dmem_n3296,
         mem_stage_inst_dmem_n3295, mem_stage_inst_dmem_n3294,
         mem_stage_inst_dmem_n3293, mem_stage_inst_dmem_n3292,
         mem_stage_inst_dmem_n3291, mem_stage_inst_dmem_n3290,
         mem_stage_inst_dmem_n3289, mem_stage_inst_dmem_n3288,
         mem_stage_inst_dmem_n3287, mem_stage_inst_dmem_n3286,
         mem_stage_inst_dmem_n3285, mem_stage_inst_dmem_n3284,
         mem_stage_inst_dmem_n3283, mem_stage_inst_dmem_n3282,
         mem_stage_inst_dmem_n3281, mem_stage_inst_dmem_n3280,
         mem_stage_inst_dmem_n3279, mem_stage_inst_dmem_n3278,
         mem_stage_inst_dmem_n3277, mem_stage_inst_dmem_n3276,
         mem_stage_inst_dmem_n3275, mem_stage_inst_dmem_n3274,
         mem_stage_inst_dmem_n3273, mem_stage_inst_dmem_n3272,
         mem_stage_inst_dmem_n3271, mem_stage_inst_dmem_n3270,
         mem_stage_inst_dmem_n3269, mem_stage_inst_dmem_n3268,
         mem_stage_inst_dmem_n3267, mem_stage_inst_dmem_n3266,
         mem_stage_inst_dmem_n3265, mem_stage_inst_dmem_n3264,
         mem_stage_inst_dmem_n3263, mem_stage_inst_dmem_n3262,
         mem_stage_inst_dmem_n3261, mem_stage_inst_dmem_n3260,
         mem_stage_inst_dmem_n3259, mem_stage_inst_dmem_n3258,
         mem_stage_inst_dmem_n3257, mem_stage_inst_dmem_n3256,
         mem_stage_inst_dmem_n3255, mem_stage_inst_dmem_n3254,
         mem_stage_inst_dmem_n3253, mem_stage_inst_dmem_n3252,
         mem_stage_inst_dmem_n3251, mem_stage_inst_dmem_n3250,
         mem_stage_inst_dmem_n3249, mem_stage_inst_dmem_n3248,
         mem_stage_inst_dmem_n3247, mem_stage_inst_dmem_n3246,
         mem_stage_inst_dmem_n3245, mem_stage_inst_dmem_n3244,
         mem_stage_inst_dmem_n3243, mem_stage_inst_dmem_n3242,
         mem_stage_inst_dmem_n3241, mem_stage_inst_dmem_n3240,
         mem_stage_inst_dmem_n3239, mem_stage_inst_dmem_n3238,
         mem_stage_inst_dmem_n3237, mem_stage_inst_dmem_n3236,
         mem_stage_inst_dmem_n3235, mem_stage_inst_dmem_n3234,
         mem_stage_inst_dmem_n3233, mem_stage_inst_dmem_n3232,
         mem_stage_inst_dmem_n3231, mem_stage_inst_dmem_n3230,
         mem_stage_inst_dmem_n3229, mem_stage_inst_dmem_n3228,
         mem_stage_inst_dmem_n3227, mem_stage_inst_dmem_n3226,
         mem_stage_inst_dmem_n3225, mem_stage_inst_dmem_n3224,
         mem_stage_inst_dmem_n3223, mem_stage_inst_dmem_n3222,
         mem_stage_inst_dmem_n3221, mem_stage_inst_dmem_n3220,
         mem_stage_inst_dmem_n3219, mem_stage_inst_dmem_n3218,
         mem_stage_inst_dmem_n3217, mem_stage_inst_dmem_n3216,
         mem_stage_inst_dmem_n3215, mem_stage_inst_dmem_n3214,
         mem_stage_inst_dmem_n3213, mem_stage_inst_dmem_n3212,
         mem_stage_inst_dmem_n3211, mem_stage_inst_dmem_n3210,
         mem_stage_inst_dmem_n3209, mem_stage_inst_dmem_n3208,
         mem_stage_inst_dmem_n3207, mem_stage_inst_dmem_n3206,
         mem_stage_inst_dmem_n3205, mem_stage_inst_dmem_n3204,
         mem_stage_inst_dmem_n3203, mem_stage_inst_dmem_n3202,
         mem_stage_inst_dmem_n3201, mem_stage_inst_dmem_n3200,
         mem_stage_inst_dmem_n3199, mem_stage_inst_dmem_n3198,
         mem_stage_inst_dmem_n3197, mem_stage_inst_dmem_n3196,
         mem_stage_inst_dmem_n3195, mem_stage_inst_dmem_n3194,
         mem_stage_inst_dmem_n3193, mem_stage_inst_dmem_n3192,
         mem_stage_inst_dmem_n3191, mem_stage_inst_dmem_n3190,
         mem_stage_inst_dmem_n3189, mem_stage_inst_dmem_n3188,
         mem_stage_inst_dmem_n3187, mem_stage_inst_dmem_n3186,
         mem_stage_inst_dmem_n3185, mem_stage_inst_dmem_n3184,
         mem_stage_inst_dmem_n3183, mem_stage_inst_dmem_n3182,
         mem_stage_inst_dmem_n3181, mem_stage_inst_dmem_n3180,
         mem_stage_inst_dmem_n3179, mem_stage_inst_dmem_n3178,
         mem_stage_inst_dmem_n3177, mem_stage_inst_dmem_n3176,
         mem_stage_inst_dmem_n3175, mem_stage_inst_dmem_n3174,
         mem_stage_inst_dmem_n3173, mem_stage_inst_dmem_n3172,
         mem_stage_inst_dmem_n3171, mem_stage_inst_dmem_n3170,
         mem_stage_inst_dmem_n3169, mem_stage_inst_dmem_n3168,
         mem_stage_inst_dmem_n3167, mem_stage_inst_dmem_n3166,
         mem_stage_inst_dmem_n3165, mem_stage_inst_dmem_n3164,
         mem_stage_inst_dmem_n3163, mem_stage_inst_dmem_n3162,
         mem_stage_inst_dmem_n3161, mem_stage_inst_dmem_n3160,
         mem_stage_inst_dmem_n3159, mem_stage_inst_dmem_n3158,
         mem_stage_inst_dmem_n3157, mem_stage_inst_dmem_n3156,
         mem_stage_inst_dmem_n3155, mem_stage_inst_dmem_n3154,
         mem_stage_inst_dmem_n3153, mem_stage_inst_dmem_n3152,
         mem_stage_inst_dmem_n3151, mem_stage_inst_dmem_n3150,
         mem_stage_inst_dmem_n3149, mem_stage_inst_dmem_n3148,
         mem_stage_inst_dmem_n3147, mem_stage_inst_dmem_n3146,
         mem_stage_inst_dmem_n3145, mem_stage_inst_dmem_n3144,
         mem_stage_inst_dmem_n3143, mem_stage_inst_dmem_n3142,
         mem_stage_inst_dmem_n3141, mem_stage_inst_dmem_n3140,
         mem_stage_inst_dmem_n3139, mem_stage_inst_dmem_n3138,
         mem_stage_inst_dmem_n3137, mem_stage_inst_dmem_n3136,
         mem_stage_inst_dmem_n3135, mem_stage_inst_dmem_n3134,
         mem_stage_inst_dmem_n3133, mem_stage_inst_dmem_n3132,
         mem_stage_inst_dmem_n3131, mem_stage_inst_dmem_n3130,
         mem_stage_inst_dmem_n3129, mem_stage_inst_dmem_n3128,
         mem_stage_inst_dmem_n3127, mem_stage_inst_dmem_n3126,
         mem_stage_inst_dmem_n3125, mem_stage_inst_dmem_n3124,
         mem_stage_inst_dmem_n3123, mem_stage_inst_dmem_n3122,
         mem_stage_inst_dmem_n3121, mem_stage_inst_dmem_n3120,
         mem_stage_inst_dmem_n3119, mem_stage_inst_dmem_n3118,
         mem_stage_inst_dmem_n3117, mem_stage_inst_dmem_n3116,
         mem_stage_inst_dmem_n3115, mem_stage_inst_dmem_n3114,
         mem_stage_inst_dmem_n3113, mem_stage_inst_dmem_n3112,
         mem_stage_inst_dmem_n3111, mem_stage_inst_dmem_n3110,
         mem_stage_inst_dmem_n3109, mem_stage_inst_dmem_n3108,
         mem_stage_inst_dmem_n3107, mem_stage_inst_dmem_n3106,
         mem_stage_inst_dmem_n3105, mem_stage_inst_dmem_n3104,
         mem_stage_inst_dmem_n3103, mem_stage_inst_dmem_n3102,
         mem_stage_inst_dmem_n3101, mem_stage_inst_dmem_n3100,
         mem_stage_inst_dmem_n3099, mem_stage_inst_dmem_n3098,
         mem_stage_inst_dmem_n3097, mem_stage_inst_dmem_n3096,
         mem_stage_inst_dmem_n3095, mem_stage_inst_dmem_n3094,
         mem_stage_inst_dmem_n3093, mem_stage_inst_dmem_n3092,
         mem_stage_inst_dmem_n3091, mem_stage_inst_dmem_n3090,
         mem_stage_inst_dmem_n3089, mem_stage_inst_dmem_n3088,
         mem_stage_inst_dmem_n3087, mem_stage_inst_dmem_n3086,
         mem_stage_inst_dmem_n3085, mem_stage_inst_dmem_n3084,
         mem_stage_inst_dmem_n3083, mem_stage_inst_dmem_n3082,
         mem_stage_inst_dmem_n3081, mem_stage_inst_dmem_n3080,
         mem_stage_inst_dmem_n3079, mem_stage_inst_dmem_n3078,
         mem_stage_inst_dmem_n3077, mem_stage_inst_dmem_n3076,
         mem_stage_inst_dmem_n3075, mem_stage_inst_dmem_n3074,
         mem_stage_inst_dmem_n3073, mem_stage_inst_dmem_n3072,
         mem_stage_inst_dmem_n3071, mem_stage_inst_dmem_n3070,
         mem_stage_inst_dmem_n3069, mem_stage_inst_dmem_n3068,
         mem_stage_inst_dmem_n3067, mem_stage_inst_dmem_n3066,
         mem_stage_inst_dmem_n3065, mem_stage_inst_dmem_n3064,
         mem_stage_inst_dmem_n3063, mem_stage_inst_dmem_n3062,
         mem_stage_inst_dmem_n3061, mem_stage_inst_dmem_n3060,
         mem_stage_inst_dmem_n3059, mem_stage_inst_dmem_n3058,
         mem_stage_inst_dmem_n3057, mem_stage_inst_dmem_n3056,
         mem_stage_inst_dmem_n3055, mem_stage_inst_dmem_n3054,
         mem_stage_inst_dmem_n3053, mem_stage_inst_dmem_n3052,
         mem_stage_inst_dmem_n3051, mem_stage_inst_dmem_n3050,
         mem_stage_inst_dmem_n3049, mem_stage_inst_dmem_n3048,
         mem_stage_inst_dmem_n3047, mem_stage_inst_dmem_n3046,
         mem_stage_inst_dmem_n3045, mem_stage_inst_dmem_n3044,
         mem_stage_inst_dmem_n3043, mem_stage_inst_dmem_n3042,
         mem_stage_inst_dmem_n3041, mem_stage_inst_dmem_n3040,
         mem_stage_inst_dmem_n3039, mem_stage_inst_dmem_n3038,
         mem_stage_inst_dmem_n3037, mem_stage_inst_dmem_n3036,
         mem_stage_inst_dmem_n3035, mem_stage_inst_dmem_n3034,
         mem_stage_inst_dmem_n3033, mem_stage_inst_dmem_n3032,
         mem_stage_inst_dmem_n3031, mem_stage_inst_dmem_n3030,
         mem_stage_inst_dmem_n3029, mem_stage_inst_dmem_n3028,
         mem_stage_inst_dmem_n3027, mem_stage_inst_dmem_n3026,
         mem_stage_inst_dmem_n3025, mem_stage_inst_dmem_n3024,
         mem_stage_inst_dmem_n3023, mem_stage_inst_dmem_n3022,
         mem_stage_inst_dmem_n3021, mem_stage_inst_dmem_n3020,
         mem_stage_inst_dmem_n3019, mem_stage_inst_dmem_n3018,
         mem_stage_inst_dmem_n3017, mem_stage_inst_dmem_n3016,
         mem_stage_inst_dmem_n3015, mem_stage_inst_dmem_n3014,
         mem_stage_inst_dmem_n3013, mem_stage_inst_dmem_n3012,
         mem_stage_inst_dmem_n3011, mem_stage_inst_dmem_n3010,
         mem_stage_inst_dmem_n3009, mem_stage_inst_dmem_n3008,
         mem_stage_inst_dmem_n3007, mem_stage_inst_dmem_n3006,
         mem_stage_inst_dmem_n3005, mem_stage_inst_dmem_n3004,
         mem_stage_inst_dmem_n3003, mem_stage_inst_dmem_n3002,
         mem_stage_inst_dmem_n3001, mem_stage_inst_dmem_n3000,
         mem_stage_inst_dmem_n2999, mem_stage_inst_dmem_n2998,
         mem_stage_inst_dmem_n2997, mem_stage_inst_dmem_n2996,
         mem_stage_inst_dmem_n2995, mem_stage_inst_dmem_n2994,
         mem_stage_inst_dmem_n2993, mem_stage_inst_dmem_n2992,
         mem_stage_inst_dmem_n2991, mem_stage_inst_dmem_n2990,
         mem_stage_inst_dmem_n2989, mem_stage_inst_dmem_n2988,
         mem_stage_inst_dmem_n2987, mem_stage_inst_dmem_n2986,
         mem_stage_inst_dmem_n2985, mem_stage_inst_dmem_n2984,
         mem_stage_inst_dmem_n2983, mem_stage_inst_dmem_n2982,
         mem_stage_inst_dmem_n2981, mem_stage_inst_dmem_n2980,
         mem_stage_inst_dmem_n2979, mem_stage_inst_dmem_n2978,
         mem_stage_inst_dmem_n2977, mem_stage_inst_dmem_n2976,
         mem_stage_inst_dmem_n2975, mem_stage_inst_dmem_n2974,
         mem_stage_inst_dmem_n2973, mem_stage_inst_dmem_n2972,
         mem_stage_inst_dmem_n2971, mem_stage_inst_dmem_n2970,
         mem_stage_inst_dmem_n2969, mem_stage_inst_dmem_n2968,
         mem_stage_inst_dmem_n2967, mem_stage_inst_dmem_n2966,
         mem_stage_inst_dmem_n2965, mem_stage_inst_dmem_n2964,
         mem_stage_inst_dmem_n2963, mem_stage_inst_dmem_n2962,
         mem_stage_inst_dmem_n2961, mem_stage_inst_dmem_n2960,
         mem_stage_inst_dmem_n2959, mem_stage_inst_dmem_n2958,
         mem_stage_inst_dmem_n2957, mem_stage_inst_dmem_n2956,
         mem_stage_inst_dmem_n2955, mem_stage_inst_dmem_n2954,
         mem_stage_inst_dmem_n2953, mem_stage_inst_dmem_n2952,
         mem_stage_inst_dmem_n2951, mem_stage_inst_dmem_n2950,
         mem_stage_inst_dmem_n2949, mem_stage_inst_dmem_n2948,
         mem_stage_inst_dmem_n2947, mem_stage_inst_dmem_n2946,
         mem_stage_inst_dmem_n2945, mem_stage_inst_dmem_n2944,
         mem_stage_inst_dmem_n2943, mem_stage_inst_dmem_n2942,
         mem_stage_inst_dmem_n2941, mem_stage_inst_dmem_n2940,
         mem_stage_inst_dmem_n2939, mem_stage_inst_dmem_n2938,
         mem_stage_inst_dmem_n2937, mem_stage_inst_dmem_n2936,
         mem_stage_inst_dmem_n2935, mem_stage_inst_dmem_n2934,
         mem_stage_inst_dmem_n2933, mem_stage_inst_dmem_n2932,
         mem_stage_inst_dmem_n2931, mem_stage_inst_dmem_n2930,
         mem_stage_inst_dmem_n2929, mem_stage_inst_dmem_n2928,
         mem_stage_inst_dmem_n2927, mem_stage_inst_dmem_n2926,
         mem_stage_inst_dmem_n2925, mem_stage_inst_dmem_n2924,
         mem_stage_inst_dmem_n2923, mem_stage_inst_dmem_n2922,
         mem_stage_inst_dmem_n2921, mem_stage_inst_dmem_n2920,
         mem_stage_inst_dmem_n2919, mem_stage_inst_dmem_n2918,
         mem_stage_inst_dmem_n2917, mem_stage_inst_dmem_n2916,
         mem_stage_inst_dmem_n2915, mem_stage_inst_dmem_n2914,
         mem_stage_inst_dmem_n2913, mem_stage_inst_dmem_n2912,
         mem_stage_inst_dmem_n2911, mem_stage_inst_dmem_n2910,
         mem_stage_inst_dmem_n2909, mem_stage_inst_dmem_n2908,
         mem_stage_inst_dmem_n2907, mem_stage_inst_dmem_n2906,
         mem_stage_inst_dmem_n2905, mem_stage_inst_dmem_n2904,
         mem_stage_inst_dmem_n2903, mem_stage_inst_dmem_n2902,
         mem_stage_inst_dmem_n2901, mem_stage_inst_dmem_n2900,
         mem_stage_inst_dmem_n2899, mem_stage_inst_dmem_n2898,
         mem_stage_inst_dmem_n2897, mem_stage_inst_dmem_n2896,
         mem_stage_inst_dmem_n2895, mem_stage_inst_dmem_n2894,
         mem_stage_inst_dmem_n2893, mem_stage_inst_dmem_n2892,
         mem_stage_inst_dmem_n2891, mem_stage_inst_dmem_n2890,
         mem_stage_inst_dmem_n2889, mem_stage_inst_dmem_n2888,
         mem_stage_inst_dmem_n2887, mem_stage_inst_dmem_n2886,
         mem_stage_inst_dmem_n2885, mem_stage_inst_dmem_n2884,
         mem_stage_inst_dmem_n2883, mem_stage_inst_dmem_n2882,
         mem_stage_inst_dmem_n2881, mem_stage_inst_dmem_n2880,
         mem_stage_inst_dmem_n2879, mem_stage_inst_dmem_n2878,
         mem_stage_inst_dmem_n2877, mem_stage_inst_dmem_n2876,
         mem_stage_inst_dmem_n2875, mem_stage_inst_dmem_n2874,
         mem_stage_inst_dmem_n2873, mem_stage_inst_dmem_n2872,
         mem_stage_inst_dmem_n2871, mem_stage_inst_dmem_n2870,
         mem_stage_inst_dmem_n2869, mem_stage_inst_dmem_n2868,
         mem_stage_inst_dmem_n2867, mem_stage_inst_dmem_n2866,
         mem_stage_inst_dmem_n2865, mem_stage_inst_dmem_n2864,
         mem_stage_inst_dmem_n2863, mem_stage_inst_dmem_n2862,
         mem_stage_inst_dmem_n2861, mem_stage_inst_dmem_n2860,
         mem_stage_inst_dmem_n2859, mem_stage_inst_dmem_n2858,
         mem_stage_inst_dmem_n2857, mem_stage_inst_dmem_n2856,
         mem_stage_inst_dmem_n2855, mem_stage_inst_dmem_n2854,
         mem_stage_inst_dmem_n2853, mem_stage_inst_dmem_n2852,
         mem_stage_inst_dmem_n2851, mem_stage_inst_dmem_n2850,
         mem_stage_inst_dmem_n2849, mem_stage_inst_dmem_n2848,
         mem_stage_inst_dmem_n2847, mem_stage_inst_dmem_n2846,
         mem_stage_inst_dmem_n2845, mem_stage_inst_dmem_n2844,
         mem_stage_inst_dmem_n2843, mem_stage_inst_dmem_n2842,
         mem_stage_inst_dmem_n2841, mem_stage_inst_dmem_n2840,
         mem_stage_inst_dmem_n2839, mem_stage_inst_dmem_n2838,
         mem_stage_inst_dmem_n2837, mem_stage_inst_dmem_n2836,
         mem_stage_inst_dmem_n2835, mem_stage_inst_dmem_n2834,
         mem_stage_inst_dmem_n2833, mem_stage_inst_dmem_n2832,
         mem_stage_inst_dmem_n2831, mem_stage_inst_dmem_n2830,
         mem_stage_inst_dmem_n2829, mem_stage_inst_dmem_n2828,
         mem_stage_inst_dmem_n2827, mem_stage_inst_dmem_n2826,
         mem_stage_inst_dmem_n2825, mem_stage_inst_dmem_n2824,
         mem_stage_inst_dmem_n2823, mem_stage_inst_dmem_n2822,
         mem_stage_inst_dmem_n2821, mem_stage_inst_dmem_n2820,
         mem_stage_inst_dmem_n2819, mem_stage_inst_dmem_n2818,
         mem_stage_inst_dmem_n2817, mem_stage_inst_dmem_n2816,
         mem_stage_inst_dmem_n2815, mem_stage_inst_dmem_n2814,
         mem_stage_inst_dmem_n2813, mem_stage_inst_dmem_n2812,
         mem_stage_inst_dmem_n2811, mem_stage_inst_dmem_n2810,
         mem_stage_inst_dmem_n2809, mem_stage_inst_dmem_n2808,
         mem_stage_inst_dmem_n2807, mem_stage_inst_dmem_n2806,
         mem_stage_inst_dmem_n2805, mem_stage_inst_dmem_n2804,
         mem_stage_inst_dmem_n2803, mem_stage_inst_dmem_n2802,
         mem_stage_inst_dmem_n2801, mem_stage_inst_dmem_n2800,
         mem_stage_inst_dmem_n2799, mem_stage_inst_dmem_n2798,
         mem_stage_inst_dmem_n2797, mem_stage_inst_dmem_n2796,
         mem_stage_inst_dmem_n2795, mem_stage_inst_dmem_n2794,
         mem_stage_inst_dmem_n2793, mem_stage_inst_dmem_n2792,
         mem_stage_inst_dmem_n2791, mem_stage_inst_dmem_n2790,
         mem_stage_inst_dmem_n2789, mem_stage_inst_dmem_n2788,
         mem_stage_inst_dmem_n2787, mem_stage_inst_dmem_n2786,
         mem_stage_inst_dmem_n2785, mem_stage_inst_dmem_n2784,
         mem_stage_inst_dmem_n2783, mem_stage_inst_dmem_n2782,
         mem_stage_inst_dmem_n2781, mem_stage_inst_dmem_n2780,
         mem_stage_inst_dmem_n2779, mem_stage_inst_dmem_n2778,
         mem_stage_inst_dmem_n2777, mem_stage_inst_dmem_n2776,
         mem_stage_inst_dmem_n2775, mem_stage_inst_dmem_n2774,
         mem_stage_inst_dmem_n2773, mem_stage_inst_dmem_n2772,
         mem_stage_inst_dmem_n2771, mem_stage_inst_dmem_n2770,
         mem_stage_inst_dmem_n2769, mem_stage_inst_dmem_n2768,
         mem_stage_inst_dmem_n2767, mem_stage_inst_dmem_n2766,
         mem_stage_inst_dmem_n2765, mem_stage_inst_dmem_n2764,
         mem_stage_inst_dmem_n2763, mem_stage_inst_dmem_n2762,
         mem_stage_inst_dmem_n2761, mem_stage_inst_dmem_n2760,
         mem_stage_inst_dmem_n2759, mem_stage_inst_dmem_n2758,
         mem_stage_inst_dmem_n2757, mem_stage_inst_dmem_n2756,
         mem_stage_inst_dmem_n2755, mem_stage_inst_dmem_n2754,
         mem_stage_inst_dmem_n2753, mem_stage_inst_dmem_n2752,
         mem_stage_inst_dmem_n2751, mem_stage_inst_dmem_n2750,
         mem_stage_inst_dmem_n2749, mem_stage_inst_dmem_n2748,
         mem_stage_inst_dmem_n2747, mem_stage_inst_dmem_n2746,
         mem_stage_inst_dmem_n2745, mem_stage_inst_dmem_n2744,
         mem_stage_inst_dmem_n2743, mem_stage_inst_dmem_n2742,
         mem_stage_inst_dmem_n2741, mem_stage_inst_dmem_n2740,
         mem_stage_inst_dmem_n2739, mem_stage_inst_dmem_n2738,
         mem_stage_inst_dmem_n2737, mem_stage_inst_dmem_n2736,
         mem_stage_inst_dmem_n2735, mem_stage_inst_dmem_n2734,
         mem_stage_inst_dmem_n2733, mem_stage_inst_dmem_n2732,
         mem_stage_inst_dmem_n2731, mem_stage_inst_dmem_n2730,
         mem_stage_inst_dmem_n2729, mem_stage_inst_dmem_n2728,
         mem_stage_inst_dmem_n2727, mem_stage_inst_dmem_n2726,
         mem_stage_inst_dmem_n2725, mem_stage_inst_dmem_n2724,
         mem_stage_inst_dmem_n2723, mem_stage_inst_dmem_n2722,
         mem_stage_inst_dmem_n2721, mem_stage_inst_dmem_n2720,
         mem_stage_inst_dmem_n2719, mem_stage_inst_dmem_n2718,
         mem_stage_inst_dmem_n2717, mem_stage_inst_dmem_n2716,
         mem_stage_inst_dmem_n2715, mem_stage_inst_dmem_n2714,
         mem_stage_inst_dmem_n2713, mem_stage_inst_dmem_n2712,
         mem_stage_inst_dmem_n2711, mem_stage_inst_dmem_n2710,
         mem_stage_inst_dmem_n2709, mem_stage_inst_dmem_n2708,
         mem_stage_inst_dmem_n2707, mem_stage_inst_dmem_n2706,
         mem_stage_inst_dmem_n2705, mem_stage_inst_dmem_n2704,
         mem_stage_inst_dmem_n2703, mem_stage_inst_dmem_n2702,
         mem_stage_inst_dmem_n2701, mem_stage_inst_dmem_n2700,
         mem_stage_inst_dmem_n2699, mem_stage_inst_dmem_n2698,
         mem_stage_inst_dmem_n2697, mem_stage_inst_dmem_n2696,
         mem_stage_inst_dmem_n2695, mem_stage_inst_dmem_n2694,
         mem_stage_inst_dmem_n2693, mem_stage_inst_dmem_n2692,
         mem_stage_inst_dmem_n2691, mem_stage_inst_dmem_n2690,
         mem_stage_inst_dmem_n2689, mem_stage_inst_dmem_n2688,
         mem_stage_inst_dmem_n2687, mem_stage_inst_dmem_n2686,
         mem_stage_inst_dmem_n2685, mem_stage_inst_dmem_n2684,
         mem_stage_inst_dmem_n2683, mem_stage_inst_dmem_n2682,
         mem_stage_inst_dmem_n2681, mem_stage_inst_dmem_n2680,
         mem_stage_inst_dmem_n2679, mem_stage_inst_dmem_n2678,
         mem_stage_inst_dmem_n2677, mem_stage_inst_dmem_n2676,
         mem_stage_inst_dmem_n2675, mem_stage_inst_dmem_n2674,
         mem_stage_inst_dmem_n2673, mem_stage_inst_dmem_n2672,
         mem_stage_inst_dmem_n2671, mem_stage_inst_dmem_n2670,
         mem_stage_inst_dmem_n2669, mem_stage_inst_dmem_n2668,
         mem_stage_inst_dmem_n2667, mem_stage_inst_dmem_n2666,
         mem_stage_inst_dmem_n2665, mem_stage_inst_dmem_n2664,
         mem_stage_inst_dmem_n2663, mem_stage_inst_dmem_n2662,
         mem_stage_inst_dmem_n2661, mem_stage_inst_dmem_n2660,
         mem_stage_inst_dmem_n2659, mem_stage_inst_dmem_n2658,
         mem_stage_inst_dmem_n2657, mem_stage_inst_dmem_n2656,
         mem_stage_inst_dmem_n2655, mem_stage_inst_dmem_n2654,
         mem_stage_inst_dmem_n2653, mem_stage_inst_dmem_n2652,
         mem_stage_inst_dmem_n2651, mem_stage_inst_dmem_n2650,
         mem_stage_inst_dmem_n2649, mem_stage_inst_dmem_n2648,
         mem_stage_inst_dmem_n2647, mem_stage_inst_dmem_n2646,
         mem_stage_inst_dmem_n2645, mem_stage_inst_dmem_n2644,
         mem_stage_inst_dmem_n2643, mem_stage_inst_dmem_n2642,
         mem_stage_inst_dmem_n2641, mem_stage_inst_dmem_n2640,
         mem_stage_inst_dmem_n2639, mem_stage_inst_dmem_n2638,
         mem_stage_inst_dmem_n2637, mem_stage_inst_dmem_n2636,
         mem_stage_inst_dmem_n2635, mem_stage_inst_dmem_n2634,
         mem_stage_inst_dmem_n2633, mem_stage_inst_dmem_n2632,
         mem_stage_inst_dmem_n2631, mem_stage_inst_dmem_n2630,
         mem_stage_inst_dmem_n2629, mem_stage_inst_dmem_n2628,
         mem_stage_inst_dmem_n2627, mem_stage_inst_dmem_n2626,
         mem_stage_inst_dmem_n2625, mem_stage_inst_dmem_n2624,
         mem_stage_inst_dmem_n2623, mem_stage_inst_dmem_n2622,
         mem_stage_inst_dmem_n2621, mem_stage_inst_dmem_n2620,
         mem_stage_inst_dmem_n2619, mem_stage_inst_dmem_n2618,
         mem_stage_inst_dmem_n2617, mem_stage_inst_dmem_n2616,
         mem_stage_inst_dmem_n2615, mem_stage_inst_dmem_n2614,
         mem_stage_inst_dmem_n2613, mem_stage_inst_dmem_n2612,
         mem_stage_inst_dmem_n2611, mem_stage_inst_dmem_n2610,
         mem_stage_inst_dmem_n2609, mem_stage_inst_dmem_n2608,
         mem_stage_inst_dmem_n2607, mem_stage_inst_dmem_n2606,
         mem_stage_inst_dmem_n2605, mem_stage_inst_dmem_n2604,
         mem_stage_inst_dmem_n2603, mem_stage_inst_dmem_n2602,
         mem_stage_inst_dmem_n2601, mem_stage_inst_dmem_n2600,
         mem_stage_inst_dmem_n2599, mem_stage_inst_dmem_n2598,
         mem_stage_inst_dmem_n2597, mem_stage_inst_dmem_n2596,
         mem_stage_inst_dmem_n2595, mem_stage_inst_dmem_n2594,
         mem_stage_inst_dmem_n2593, mem_stage_inst_dmem_n2592,
         mem_stage_inst_dmem_n2591, mem_stage_inst_dmem_n2590,
         mem_stage_inst_dmem_n2589, mem_stage_inst_dmem_n2588,
         mem_stage_inst_dmem_n2587, mem_stage_inst_dmem_n2586,
         mem_stage_inst_dmem_n2585, mem_stage_inst_dmem_n2584,
         mem_stage_inst_dmem_n2583, mem_stage_inst_dmem_n2582,
         mem_stage_inst_dmem_n2581, mem_stage_inst_dmem_n2580,
         mem_stage_inst_dmem_n2579, mem_stage_inst_dmem_n2578,
         mem_stage_inst_dmem_n2577, mem_stage_inst_dmem_n2576,
         mem_stage_inst_dmem_n2575, mem_stage_inst_dmem_n2574,
         mem_stage_inst_dmem_n2573, mem_stage_inst_dmem_n2572,
         mem_stage_inst_dmem_n2571, mem_stage_inst_dmem_n2570,
         mem_stage_inst_dmem_n2569, mem_stage_inst_dmem_n2568,
         mem_stage_inst_dmem_n2567, mem_stage_inst_dmem_n2566,
         mem_stage_inst_dmem_n2565, mem_stage_inst_dmem_n2564,
         mem_stage_inst_dmem_n2563, mem_stage_inst_dmem_n2562,
         mem_stage_inst_dmem_n2561, mem_stage_inst_dmem_n2560,
         mem_stage_inst_dmem_n2559, mem_stage_inst_dmem_n2558,
         mem_stage_inst_dmem_n2557, mem_stage_inst_dmem_n2556,
         mem_stage_inst_dmem_n2555, mem_stage_inst_dmem_n2554,
         mem_stage_inst_dmem_n2553, mem_stage_inst_dmem_n2552,
         mem_stage_inst_dmem_n2551, mem_stage_inst_dmem_n2550,
         mem_stage_inst_dmem_n2549, mem_stage_inst_dmem_n2548,
         mem_stage_inst_dmem_n2547, mem_stage_inst_dmem_n2546,
         mem_stage_inst_dmem_n2545, mem_stage_inst_dmem_n2544,
         mem_stage_inst_dmem_n2543, mem_stage_inst_dmem_n2542,
         mem_stage_inst_dmem_n2541, mem_stage_inst_dmem_n2540,
         mem_stage_inst_dmem_n2539, mem_stage_inst_dmem_n2538,
         mem_stage_inst_dmem_n2537, mem_stage_inst_dmem_n2536,
         mem_stage_inst_dmem_n2535, mem_stage_inst_dmem_n2534,
         mem_stage_inst_dmem_n2533, mem_stage_inst_dmem_n2532,
         mem_stage_inst_dmem_n2531, mem_stage_inst_dmem_n2530,
         mem_stage_inst_dmem_n2529, mem_stage_inst_dmem_n2528,
         mem_stage_inst_dmem_n2527, mem_stage_inst_dmem_n2526,
         mem_stage_inst_dmem_n2525, mem_stage_inst_dmem_n2524,
         mem_stage_inst_dmem_n2523, mem_stage_inst_dmem_n2522,
         mem_stage_inst_dmem_n2521, mem_stage_inst_dmem_n2520,
         mem_stage_inst_dmem_n2519, mem_stage_inst_dmem_n2518,
         mem_stage_inst_dmem_n2517, mem_stage_inst_dmem_n2516,
         mem_stage_inst_dmem_n2515, mem_stage_inst_dmem_n2514,
         mem_stage_inst_dmem_n2513, mem_stage_inst_dmem_n2512,
         mem_stage_inst_dmem_n2511, mem_stage_inst_dmem_n2510,
         mem_stage_inst_dmem_n2509, mem_stage_inst_dmem_n2508,
         mem_stage_inst_dmem_n2507, mem_stage_inst_dmem_n2506,
         mem_stage_inst_dmem_n2505, mem_stage_inst_dmem_n2504,
         mem_stage_inst_dmem_n2503, mem_stage_inst_dmem_n2502,
         mem_stage_inst_dmem_n2501, mem_stage_inst_dmem_n2500,
         mem_stage_inst_dmem_n2499, mem_stage_inst_dmem_n2498,
         mem_stage_inst_dmem_n2497, mem_stage_inst_dmem_n2496,
         mem_stage_inst_dmem_n2495, mem_stage_inst_dmem_n2494,
         mem_stage_inst_dmem_n2493, mem_stage_inst_dmem_n2492,
         mem_stage_inst_dmem_n2491, mem_stage_inst_dmem_n2490,
         mem_stage_inst_dmem_n2489, mem_stage_inst_dmem_n2488,
         mem_stage_inst_dmem_n2487, mem_stage_inst_dmem_n2486,
         mem_stage_inst_dmem_n2485, mem_stage_inst_dmem_n2484,
         mem_stage_inst_dmem_n2483, mem_stage_inst_dmem_n2482,
         mem_stage_inst_dmem_n2481, mem_stage_inst_dmem_n2480,
         mem_stage_inst_dmem_n2479, mem_stage_inst_dmem_n2478,
         mem_stage_inst_dmem_n2477, mem_stage_inst_dmem_n2476,
         mem_stage_inst_dmem_n2475, mem_stage_inst_dmem_n2474,
         mem_stage_inst_dmem_n2473, mem_stage_inst_dmem_n2472,
         mem_stage_inst_dmem_n2471, mem_stage_inst_dmem_n2470,
         mem_stage_inst_dmem_n2469, mem_stage_inst_dmem_n2468,
         mem_stage_inst_dmem_n2467, mem_stage_inst_dmem_n2466,
         mem_stage_inst_dmem_n2465, mem_stage_inst_dmem_n2464,
         mem_stage_inst_dmem_n2463, mem_stage_inst_dmem_n2462,
         mem_stage_inst_dmem_n2461, mem_stage_inst_dmem_n2460,
         mem_stage_inst_dmem_n2459, mem_stage_inst_dmem_n2458,
         mem_stage_inst_dmem_n2457, mem_stage_inst_dmem_n2456,
         mem_stage_inst_dmem_n2455, mem_stage_inst_dmem_n2454,
         mem_stage_inst_dmem_n2453, mem_stage_inst_dmem_n2452,
         mem_stage_inst_dmem_n2451, mem_stage_inst_dmem_n2450,
         mem_stage_inst_dmem_n2449, mem_stage_inst_dmem_n2448,
         mem_stage_inst_dmem_n2447, mem_stage_inst_dmem_n2446,
         mem_stage_inst_dmem_n2445, mem_stage_inst_dmem_n2444,
         mem_stage_inst_dmem_n2443, mem_stage_inst_dmem_n2442,
         mem_stage_inst_dmem_n2441, mem_stage_inst_dmem_n2440,
         mem_stage_inst_dmem_n2439, mem_stage_inst_dmem_n2438,
         mem_stage_inst_dmem_n2437, mem_stage_inst_dmem_n2436,
         mem_stage_inst_dmem_n2435, mem_stage_inst_dmem_n2434,
         mem_stage_inst_dmem_n2433, mem_stage_inst_dmem_n2432,
         mem_stage_inst_dmem_n2431, mem_stage_inst_dmem_n2430,
         mem_stage_inst_dmem_n2429, mem_stage_inst_dmem_n2428,
         mem_stage_inst_dmem_n2427, mem_stage_inst_dmem_n2426,
         mem_stage_inst_dmem_n2425, mem_stage_inst_dmem_n2424,
         mem_stage_inst_dmem_n2423, mem_stage_inst_dmem_n2422,
         mem_stage_inst_dmem_n2421, mem_stage_inst_dmem_n2420,
         mem_stage_inst_dmem_n2419, mem_stage_inst_dmem_n2418,
         mem_stage_inst_dmem_n2417, mem_stage_inst_dmem_n2416,
         mem_stage_inst_dmem_n2415, mem_stage_inst_dmem_n2414,
         mem_stage_inst_dmem_n2413, mem_stage_inst_dmem_n2412,
         mem_stage_inst_dmem_n2411, mem_stage_inst_dmem_n2410,
         mem_stage_inst_dmem_n2409, mem_stage_inst_dmem_n2408,
         mem_stage_inst_dmem_n2407, mem_stage_inst_dmem_n2406,
         mem_stage_inst_dmem_n2405, mem_stage_inst_dmem_n2404,
         mem_stage_inst_dmem_n2403, mem_stage_inst_dmem_n2402,
         mem_stage_inst_dmem_n2401, mem_stage_inst_dmem_n2400,
         mem_stage_inst_dmem_n2399, mem_stage_inst_dmem_n2398,
         mem_stage_inst_dmem_n2397, mem_stage_inst_dmem_n2396,
         mem_stage_inst_dmem_n2395, mem_stage_inst_dmem_n2394,
         mem_stage_inst_dmem_n2393, mem_stage_inst_dmem_n2392,
         mem_stage_inst_dmem_n2391, mem_stage_inst_dmem_n2390,
         mem_stage_inst_dmem_n2389, mem_stage_inst_dmem_n2388,
         mem_stage_inst_dmem_n2387, mem_stage_inst_dmem_n2386,
         mem_stage_inst_dmem_n2385, mem_stage_inst_dmem_n2384,
         mem_stage_inst_dmem_n2383, mem_stage_inst_dmem_n2382,
         mem_stage_inst_dmem_n2381, mem_stage_inst_dmem_n2380,
         mem_stage_inst_dmem_n2379, mem_stage_inst_dmem_n2378,
         mem_stage_inst_dmem_n2377, mem_stage_inst_dmem_n2376,
         mem_stage_inst_dmem_n2375, mem_stage_inst_dmem_n2374,
         mem_stage_inst_dmem_n2373, mem_stage_inst_dmem_n2372,
         mem_stage_inst_dmem_n2371, mem_stage_inst_dmem_n2370,
         mem_stage_inst_dmem_n2369, mem_stage_inst_dmem_n2368,
         mem_stage_inst_dmem_n2367, mem_stage_inst_dmem_n2366,
         mem_stage_inst_dmem_n2365, mem_stage_inst_dmem_n2364,
         mem_stage_inst_dmem_n2363, mem_stage_inst_dmem_n2362,
         mem_stage_inst_dmem_n2361, mem_stage_inst_dmem_n2360,
         mem_stage_inst_dmem_n2359, mem_stage_inst_dmem_n2358,
         mem_stage_inst_dmem_n2357, mem_stage_inst_dmem_n2356,
         mem_stage_inst_dmem_n2355, mem_stage_inst_dmem_n2354,
         mem_stage_inst_dmem_n2353, mem_stage_inst_dmem_n2352,
         mem_stage_inst_dmem_n2351, mem_stage_inst_dmem_n2350,
         mem_stage_inst_dmem_n2349, mem_stage_inst_dmem_n2348,
         mem_stage_inst_dmem_n2347, mem_stage_inst_dmem_n2346,
         mem_stage_inst_dmem_n2345, mem_stage_inst_dmem_n2344,
         mem_stage_inst_dmem_n2343, mem_stage_inst_dmem_n2342,
         mem_stage_inst_dmem_n2341, mem_stage_inst_dmem_n2340,
         mem_stage_inst_dmem_n2339, mem_stage_inst_dmem_n2338,
         mem_stage_inst_dmem_n2337, mem_stage_inst_dmem_n2336,
         mem_stage_inst_dmem_n2335, mem_stage_inst_dmem_n2334,
         mem_stage_inst_dmem_n2333, mem_stage_inst_dmem_n2332,
         mem_stage_inst_dmem_n2331, mem_stage_inst_dmem_n2330,
         mem_stage_inst_dmem_n2329, mem_stage_inst_dmem_n2328,
         mem_stage_inst_dmem_n2327, mem_stage_inst_dmem_n2326,
         mem_stage_inst_dmem_n2325, mem_stage_inst_dmem_n2324,
         mem_stage_inst_dmem_n2323, mem_stage_inst_dmem_n2322,
         mem_stage_inst_dmem_n2321, mem_stage_inst_dmem_n2320,
         mem_stage_inst_dmem_n2319, mem_stage_inst_dmem_n2318,
         mem_stage_inst_dmem_n2317, mem_stage_inst_dmem_n2316,
         mem_stage_inst_dmem_n2315, mem_stage_inst_dmem_n2314,
         mem_stage_inst_dmem_n2313, mem_stage_inst_dmem_n2312,
         mem_stage_inst_dmem_n2311, mem_stage_inst_dmem_n2310,
         mem_stage_inst_dmem_n2309, mem_stage_inst_dmem_n2308,
         mem_stage_inst_dmem_n2307, mem_stage_inst_dmem_n2306,
         mem_stage_inst_dmem_n2305, mem_stage_inst_dmem_n2304,
         mem_stage_inst_dmem_n2303, mem_stage_inst_dmem_n2302,
         mem_stage_inst_dmem_n2301, mem_stage_inst_dmem_n2300,
         mem_stage_inst_dmem_n2299, mem_stage_inst_dmem_n2298,
         mem_stage_inst_dmem_n2297, mem_stage_inst_dmem_n2296,
         mem_stage_inst_dmem_n2295, mem_stage_inst_dmem_n2294,
         mem_stage_inst_dmem_n2293, mem_stage_inst_dmem_n2292,
         mem_stage_inst_dmem_n2291, mem_stage_inst_dmem_n2290,
         mem_stage_inst_dmem_n2289, mem_stage_inst_dmem_n2288,
         mem_stage_inst_dmem_n2287, mem_stage_inst_dmem_n2286,
         mem_stage_inst_dmem_n2285, mem_stage_inst_dmem_n2284,
         mem_stage_inst_dmem_n2283, mem_stage_inst_dmem_n2282,
         mem_stage_inst_dmem_n2281, mem_stage_inst_dmem_n2280,
         mem_stage_inst_dmem_n2279, mem_stage_inst_dmem_n2278,
         mem_stage_inst_dmem_n2277, mem_stage_inst_dmem_n2276,
         mem_stage_inst_dmem_n2275, mem_stage_inst_dmem_n2274,
         mem_stage_inst_dmem_n2273, mem_stage_inst_dmem_n2272,
         mem_stage_inst_dmem_n2271, mem_stage_inst_dmem_n2270,
         mem_stage_inst_dmem_n2269, mem_stage_inst_dmem_n2268,
         mem_stage_inst_dmem_n2267, mem_stage_inst_dmem_n2266,
         mem_stage_inst_dmem_n2265, mem_stage_inst_dmem_n2264,
         mem_stage_inst_dmem_n2263, mem_stage_inst_dmem_n2262,
         mem_stage_inst_dmem_n2261, mem_stage_inst_dmem_n2260,
         mem_stage_inst_dmem_n2259, mem_stage_inst_dmem_n2258,
         mem_stage_inst_dmem_n2257, mem_stage_inst_dmem_n2256,
         mem_stage_inst_dmem_n2255, mem_stage_inst_dmem_n2254,
         mem_stage_inst_dmem_n2253, mem_stage_inst_dmem_n2252,
         mem_stage_inst_dmem_n2251, mem_stage_inst_dmem_n2250,
         mem_stage_inst_dmem_n2249, mem_stage_inst_dmem_n2248,
         mem_stage_inst_dmem_n2247, mem_stage_inst_dmem_n2246,
         mem_stage_inst_dmem_n2245, mem_stage_inst_dmem_n2244,
         mem_stage_inst_dmem_n2243, mem_stage_inst_dmem_n2242,
         mem_stage_inst_dmem_n2241, mem_stage_inst_dmem_n2240,
         mem_stage_inst_dmem_n2239, mem_stage_inst_dmem_n2238,
         mem_stage_inst_dmem_n2237, mem_stage_inst_dmem_n2236,
         mem_stage_inst_dmem_n2235, mem_stage_inst_dmem_n2234,
         mem_stage_inst_dmem_n2233, mem_stage_inst_dmem_n2232,
         mem_stage_inst_dmem_n2231, mem_stage_inst_dmem_n2230,
         mem_stage_inst_dmem_n2229, mem_stage_inst_dmem_n2228,
         mem_stage_inst_dmem_n2227, mem_stage_inst_dmem_n2226,
         mem_stage_inst_dmem_n2225, mem_stage_inst_dmem_n2224,
         mem_stage_inst_dmem_n2223, mem_stage_inst_dmem_n2222,
         mem_stage_inst_dmem_n2221, mem_stage_inst_dmem_n2220,
         mem_stage_inst_dmem_n2219, mem_stage_inst_dmem_n2218,
         mem_stage_inst_dmem_n2217, mem_stage_inst_dmem_n2216,
         mem_stage_inst_dmem_n2215, mem_stage_inst_dmem_n2214,
         mem_stage_inst_dmem_n2213, mem_stage_inst_dmem_n2212,
         mem_stage_inst_dmem_n2211, mem_stage_inst_dmem_n2210,
         mem_stage_inst_dmem_n2209, mem_stage_inst_dmem_n2208,
         mem_stage_inst_dmem_n2207, mem_stage_inst_dmem_n2206,
         mem_stage_inst_dmem_n2205, mem_stage_inst_dmem_n2204,
         mem_stage_inst_dmem_n2203, mem_stage_inst_dmem_n2202,
         mem_stage_inst_dmem_n2201, mem_stage_inst_dmem_n2200,
         mem_stage_inst_dmem_n2199, mem_stage_inst_dmem_n2198,
         mem_stage_inst_dmem_n2197, mem_stage_inst_dmem_n2196,
         mem_stage_inst_dmem_n2195, mem_stage_inst_dmem_n2194,
         mem_stage_inst_dmem_n2193, mem_stage_inst_dmem_n2192,
         mem_stage_inst_dmem_n2191, mem_stage_inst_dmem_n2190,
         mem_stage_inst_dmem_n2189, mem_stage_inst_dmem_n2188,
         mem_stage_inst_dmem_n2187, mem_stage_inst_dmem_n2186,
         mem_stage_inst_dmem_n2185, mem_stage_inst_dmem_n2184,
         mem_stage_inst_dmem_n2183, mem_stage_inst_dmem_n2182,
         mem_stage_inst_dmem_n2181, mem_stage_inst_dmem_n2180,
         mem_stage_inst_dmem_n2179, mem_stage_inst_dmem_n2178,
         mem_stage_inst_dmem_n2177, mem_stage_inst_dmem_n2176,
         mem_stage_inst_dmem_n2175, mem_stage_inst_dmem_n2174,
         mem_stage_inst_dmem_n2173, mem_stage_inst_dmem_n2172,
         mem_stage_inst_dmem_n2171, mem_stage_inst_dmem_n2170,
         mem_stage_inst_dmem_n2169, mem_stage_inst_dmem_n2168,
         mem_stage_inst_dmem_n2167, mem_stage_inst_dmem_n2166,
         mem_stage_inst_dmem_n2165, mem_stage_inst_dmem_n2164,
         mem_stage_inst_dmem_n2163, mem_stage_inst_dmem_n2162,
         mem_stage_inst_dmem_n2161, mem_stage_inst_dmem_n2160,
         mem_stage_inst_dmem_n2159, mem_stage_inst_dmem_n2158,
         mem_stage_inst_dmem_n2157, mem_stage_inst_dmem_n2156,
         mem_stage_inst_dmem_n2155, mem_stage_inst_dmem_n2154,
         mem_stage_inst_dmem_n2153, mem_stage_inst_dmem_n2152,
         mem_stage_inst_dmem_n2151, mem_stage_inst_dmem_n2150,
         mem_stage_inst_dmem_n2149, mem_stage_inst_dmem_n2148,
         mem_stage_inst_dmem_n2147, mem_stage_inst_dmem_n2146,
         mem_stage_inst_dmem_n2145, mem_stage_inst_dmem_n2144,
         mem_stage_inst_dmem_n2143, mem_stage_inst_dmem_n2142,
         mem_stage_inst_dmem_n2141, mem_stage_inst_dmem_n2140,
         mem_stage_inst_dmem_n2139, mem_stage_inst_dmem_n2138,
         mem_stage_inst_dmem_n2137, mem_stage_inst_dmem_n2136,
         mem_stage_inst_dmem_n2135, mem_stage_inst_dmem_n2134,
         mem_stage_inst_dmem_n2133, mem_stage_inst_dmem_n2132,
         mem_stage_inst_dmem_n2131, mem_stage_inst_dmem_n2130,
         mem_stage_inst_dmem_n2129, mem_stage_inst_dmem_n2128,
         mem_stage_inst_dmem_n2127, mem_stage_inst_dmem_n2126,
         mem_stage_inst_dmem_n2125, mem_stage_inst_dmem_n2124,
         mem_stage_inst_dmem_n2123, mem_stage_inst_dmem_n2122,
         mem_stage_inst_dmem_n2121, mem_stage_inst_dmem_n2120,
         mem_stage_inst_dmem_n2119, mem_stage_inst_dmem_n2118,
         mem_stage_inst_dmem_n2117, mem_stage_inst_dmem_n2116,
         mem_stage_inst_dmem_n2115, mem_stage_inst_dmem_n2114,
         mem_stage_inst_dmem_n2113, mem_stage_inst_dmem_n2112,
         mem_stage_inst_dmem_n2111, mem_stage_inst_dmem_n2110,
         mem_stage_inst_dmem_n2109, mem_stage_inst_dmem_n2108,
         mem_stage_inst_dmem_n2107, mem_stage_inst_dmem_n2106,
         mem_stage_inst_dmem_n2105, mem_stage_inst_dmem_n2104,
         mem_stage_inst_dmem_n2103, mem_stage_inst_dmem_n2102,
         mem_stage_inst_dmem_n2101, mem_stage_inst_dmem_n2100,
         mem_stage_inst_dmem_n2099, mem_stage_inst_dmem_n2098,
         mem_stage_inst_dmem_n2097, mem_stage_inst_dmem_n2096,
         mem_stage_inst_dmem_n2095, mem_stage_inst_dmem_n2094,
         mem_stage_inst_dmem_n2093, mem_stage_inst_dmem_n2092,
         mem_stage_inst_dmem_n2091, mem_stage_inst_dmem_n2090,
         mem_stage_inst_dmem_n2089, mem_stage_inst_dmem_n2088,
         mem_stage_inst_dmem_n2087, mem_stage_inst_dmem_n2086,
         mem_stage_inst_dmem_n2085, mem_stage_inst_dmem_n2084,
         mem_stage_inst_dmem_n2083, mem_stage_inst_dmem_n2082,
         mem_stage_inst_dmem_n2081, mem_stage_inst_dmem_n2080,
         mem_stage_inst_dmem_n2079, mem_stage_inst_dmem_n2078,
         mem_stage_inst_dmem_n2077, mem_stage_inst_dmem_n2076,
         mem_stage_inst_dmem_n2075, mem_stage_inst_dmem_n2074,
         mem_stage_inst_dmem_n2073, mem_stage_inst_dmem_n2072,
         mem_stage_inst_dmem_n2071, mem_stage_inst_dmem_n2070,
         mem_stage_inst_dmem_n2069, mem_stage_inst_dmem_n2068,
         mem_stage_inst_dmem_n2067, mem_stage_inst_dmem_n2066,
         mem_stage_inst_dmem_n2065, mem_stage_inst_dmem_n2064,
         mem_stage_inst_dmem_n2063, mem_stage_inst_dmem_n2062,
         mem_stage_inst_dmem_n2061, mem_stage_inst_dmem_n2060,
         mem_stage_inst_dmem_n2059, mem_stage_inst_dmem_n2058,
         mem_stage_inst_dmem_n2057, mem_stage_inst_dmem_n2056,
         mem_stage_inst_dmem_n2055, mem_stage_inst_dmem_n2054,
         mem_stage_inst_dmem_n2053, mem_stage_inst_dmem_n2052,
         mem_stage_inst_dmem_n2051, mem_stage_inst_dmem_n2050,
         mem_stage_inst_dmem_n2049, mem_stage_inst_dmem_n2048,
         mem_stage_inst_dmem_n2047, mem_stage_inst_dmem_n2046,
         mem_stage_inst_dmem_n2045, mem_stage_inst_dmem_n2044,
         mem_stage_inst_dmem_n2043, mem_stage_inst_dmem_n2042,
         mem_stage_inst_dmem_n2041, mem_stage_inst_dmem_n2040,
         mem_stage_inst_dmem_n2039, mem_stage_inst_dmem_n2038,
         mem_stage_inst_dmem_n2037, mem_stage_inst_dmem_n2036,
         mem_stage_inst_dmem_n2035, mem_stage_inst_dmem_n2034,
         mem_stage_inst_dmem_n2033, mem_stage_inst_dmem_n2032,
         mem_stage_inst_dmem_n2031, mem_stage_inst_dmem_n2030,
         mem_stage_inst_dmem_n2029, mem_stage_inst_dmem_n2028,
         mem_stage_inst_dmem_n2027, mem_stage_inst_dmem_n2026,
         mem_stage_inst_dmem_n2025, mem_stage_inst_dmem_n2024,
         mem_stage_inst_dmem_n2023, mem_stage_inst_dmem_n2022,
         mem_stage_inst_dmem_n2021, mem_stage_inst_dmem_n2020,
         mem_stage_inst_dmem_n2019, mem_stage_inst_dmem_n2018,
         mem_stage_inst_dmem_n2017, mem_stage_inst_dmem_n2016,
         mem_stage_inst_dmem_n2015, mem_stage_inst_dmem_n2014,
         mem_stage_inst_dmem_n2013, mem_stage_inst_dmem_n2012,
         mem_stage_inst_dmem_n2011, mem_stage_inst_dmem_n2010,
         mem_stage_inst_dmem_n2009, mem_stage_inst_dmem_n2008,
         mem_stage_inst_dmem_n2007, mem_stage_inst_dmem_n2006,
         mem_stage_inst_dmem_n2005, mem_stage_inst_dmem_n2004,
         mem_stage_inst_dmem_n2003, mem_stage_inst_dmem_n2002,
         mem_stage_inst_dmem_n2001, mem_stage_inst_dmem_n2000,
         mem_stage_inst_dmem_n1999, mem_stage_inst_dmem_n1998,
         mem_stage_inst_dmem_n1997, mem_stage_inst_dmem_n1996,
         mem_stage_inst_dmem_n1995, mem_stage_inst_dmem_n1994,
         mem_stage_inst_dmem_n1993, mem_stage_inst_dmem_n1992,
         mem_stage_inst_dmem_n1991, mem_stage_inst_dmem_n1990,
         mem_stage_inst_dmem_n1989, mem_stage_inst_dmem_n1988,
         mem_stage_inst_dmem_n1987, mem_stage_inst_dmem_n1986,
         mem_stage_inst_dmem_n1985, mem_stage_inst_dmem_n1984,
         mem_stage_inst_dmem_n1983, mem_stage_inst_dmem_n1982,
         mem_stage_inst_dmem_n1981, mem_stage_inst_dmem_n1980,
         mem_stage_inst_dmem_n1979, mem_stage_inst_dmem_n1978,
         mem_stage_inst_dmem_n1977, mem_stage_inst_dmem_n1976,
         mem_stage_inst_dmem_n1975, mem_stage_inst_dmem_n1974,
         mem_stage_inst_dmem_n1973, mem_stage_inst_dmem_n1972,
         mem_stage_inst_dmem_n1971, mem_stage_inst_dmem_n1970,
         mem_stage_inst_dmem_n1969, mem_stage_inst_dmem_n1968,
         mem_stage_inst_dmem_n1967, mem_stage_inst_dmem_n1966,
         mem_stage_inst_dmem_n1965, mem_stage_inst_dmem_n1964,
         mem_stage_inst_dmem_n1963, mem_stage_inst_dmem_n1962,
         mem_stage_inst_dmem_n1961, mem_stage_inst_dmem_n1960,
         mem_stage_inst_dmem_n1959, mem_stage_inst_dmem_n1958,
         mem_stage_inst_dmem_n1957, mem_stage_inst_dmem_n1956,
         mem_stage_inst_dmem_n1955, mem_stage_inst_dmem_n1954,
         mem_stage_inst_dmem_n1953, mem_stage_inst_dmem_n1952,
         mem_stage_inst_dmem_n1951, mem_stage_inst_dmem_n1950,
         mem_stage_inst_dmem_n1949, mem_stage_inst_dmem_n1948,
         mem_stage_inst_dmem_n1947, mem_stage_inst_dmem_n1946,
         mem_stage_inst_dmem_n1945, mem_stage_inst_dmem_n1944,
         mem_stage_inst_dmem_n1943, mem_stage_inst_dmem_n1942,
         mem_stage_inst_dmem_n1941, mem_stage_inst_dmem_n1940,
         mem_stage_inst_dmem_n1939, mem_stage_inst_dmem_n1938,
         mem_stage_inst_dmem_n1937, mem_stage_inst_dmem_n1936,
         mem_stage_inst_dmem_n1935, mem_stage_inst_dmem_n1934,
         mem_stage_inst_dmem_n1933, mem_stage_inst_dmem_n1932,
         mem_stage_inst_dmem_n1931, mem_stage_inst_dmem_n1930,
         mem_stage_inst_dmem_n1929, mem_stage_inst_dmem_n1928,
         mem_stage_inst_dmem_n1927, mem_stage_inst_dmem_n1926,
         mem_stage_inst_dmem_n1925, mem_stage_inst_dmem_n1924,
         mem_stage_inst_dmem_n1923, mem_stage_inst_dmem_n1922,
         mem_stage_inst_dmem_n1921, mem_stage_inst_dmem_n1920,
         mem_stage_inst_dmem_n1919, mem_stage_inst_dmem_n1918,
         mem_stage_inst_dmem_n1917, mem_stage_inst_dmem_n1916,
         mem_stage_inst_dmem_n1915, mem_stage_inst_dmem_n1914,
         mem_stage_inst_dmem_n1913, mem_stage_inst_dmem_n1912,
         mem_stage_inst_dmem_n1911, mem_stage_inst_dmem_n1910,
         mem_stage_inst_dmem_n1909, mem_stage_inst_dmem_n1908,
         mem_stage_inst_dmem_n1907, mem_stage_inst_dmem_n1906,
         mem_stage_inst_dmem_n1905, mem_stage_inst_dmem_n1904,
         mem_stage_inst_dmem_n1903, mem_stage_inst_dmem_n1902,
         mem_stage_inst_dmem_n1901, mem_stage_inst_dmem_n1900,
         mem_stage_inst_dmem_n1899, mem_stage_inst_dmem_n1898,
         mem_stage_inst_dmem_n1897, mem_stage_inst_dmem_n1896,
         mem_stage_inst_dmem_n1895, mem_stage_inst_dmem_n1894,
         mem_stage_inst_dmem_n1893, mem_stage_inst_dmem_n1892,
         mem_stage_inst_dmem_n1891, mem_stage_inst_dmem_n1890,
         mem_stage_inst_dmem_n1889, mem_stage_inst_dmem_n1888,
         mem_stage_inst_dmem_n1887, mem_stage_inst_dmem_n1886,
         mem_stage_inst_dmem_n1885, mem_stage_inst_dmem_n1884,
         mem_stage_inst_dmem_n1883, mem_stage_inst_dmem_n1882,
         mem_stage_inst_dmem_n1881, mem_stage_inst_dmem_n1880,
         mem_stage_inst_dmem_n1879, mem_stage_inst_dmem_n1878,
         mem_stage_inst_dmem_n1877, mem_stage_inst_dmem_n1876,
         mem_stage_inst_dmem_n1875, mem_stage_inst_dmem_n1874,
         mem_stage_inst_dmem_n1873, mem_stage_inst_dmem_n1872,
         mem_stage_inst_dmem_n1871, mem_stage_inst_dmem_n1870,
         mem_stage_inst_dmem_n1869, mem_stage_inst_dmem_n1868,
         mem_stage_inst_dmem_n1867, mem_stage_inst_dmem_n1866,
         mem_stage_inst_dmem_n1865, mem_stage_inst_dmem_n1864,
         mem_stage_inst_dmem_n1863, mem_stage_inst_dmem_n1862,
         mem_stage_inst_dmem_n1861, mem_stage_inst_dmem_n1860,
         mem_stage_inst_dmem_n1859, mem_stage_inst_dmem_n1858,
         mem_stage_inst_dmem_n1857, mem_stage_inst_dmem_n1856,
         mem_stage_inst_dmem_n1855, mem_stage_inst_dmem_n1854,
         mem_stage_inst_dmem_n1853, mem_stage_inst_dmem_n1852,
         mem_stage_inst_dmem_n1851, mem_stage_inst_dmem_n1850,
         mem_stage_inst_dmem_n1849, mem_stage_inst_dmem_n1848,
         mem_stage_inst_dmem_n1847, mem_stage_inst_dmem_n1846,
         mem_stage_inst_dmem_n1845, mem_stage_inst_dmem_n1844,
         mem_stage_inst_dmem_n1843, mem_stage_inst_dmem_n1842,
         mem_stage_inst_dmem_n1841, mem_stage_inst_dmem_n1840,
         mem_stage_inst_dmem_n1839, mem_stage_inst_dmem_n1838,
         mem_stage_inst_dmem_n1837, mem_stage_inst_dmem_n1836,
         mem_stage_inst_dmem_n1835, mem_stage_inst_dmem_n1834,
         mem_stage_inst_dmem_n1833, mem_stage_inst_dmem_n1832,
         mem_stage_inst_dmem_n1831, mem_stage_inst_dmem_n1830,
         mem_stage_inst_dmem_n1829, mem_stage_inst_dmem_n1828,
         mem_stage_inst_dmem_n1827, mem_stage_inst_dmem_n1826,
         mem_stage_inst_dmem_n1825, mem_stage_inst_dmem_n1824,
         mem_stage_inst_dmem_n1823, mem_stage_inst_dmem_n1822,
         mem_stage_inst_dmem_n1821, mem_stage_inst_dmem_n1820,
         mem_stage_inst_dmem_n1819, mem_stage_inst_dmem_n1818,
         mem_stage_inst_dmem_n1817, mem_stage_inst_dmem_n1816,
         mem_stage_inst_dmem_n1815, mem_stage_inst_dmem_n1814,
         mem_stage_inst_dmem_n1813, mem_stage_inst_dmem_n1812,
         mem_stage_inst_dmem_n1811, mem_stage_inst_dmem_n1810,
         mem_stage_inst_dmem_n1809, mem_stage_inst_dmem_n1808,
         mem_stage_inst_dmem_n1807, mem_stage_inst_dmem_n1806,
         mem_stage_inst_dmem_n1805, mem_stage_inst_dmem_n1804,
         mem_stage_inst_dmem_n1803, mem_stage_inst_dmem_n1802,
         mem_stage_inst_dmem_n1801, mem_stage_inst_dmem_n1800,
         mem_stage_inst_dmem_n1799, mem_stage_inst_dmem_n1798,
         mem_stage_inst_dmem_n1797, mem_stage_inst_dmem_n1796,
         mem_stage_inst_dmem_n1795, mem_stage_inst_dmem_n1794,
         mem_stage_inst_dmem_n1793, mem_stage_inst_dmem_n1792,
         mem_stage_inst_dmem_n1791, mem_stage_inst_dmem_n1790,
         mem_stage_inst_dmem_n1789, mem_stage_inst_dmem_n1788,
         mem_stage_inst_dmem_n1787, mem_stage_inst_dmem_n1786,
         mem_stage_inst_dmem_n1785, mem_stage_inst_dmem_n1784,
         mem_stage_inst_dmem_n1783, mem_stage_inst_dmem_n1782,
         mem_stage_inst_dmem_n1781, mem_stage_inst_dmem_n1780,
         mem_stage_inst_dmem_n1779, mem_stage_inst_dmem_n1778,
         mem_stage_inst_dmem_n1777, mem_stage_inst_dmem_n1776,
         mem_stage_inst_dmem_n1775, mem_stage_inst_dmem_n1774,
         mem_stage_inst_dmem_n1773, mem_stage_inst_dmem_n1772,
         mem_stage_inst_dmem_n1771, mem_stage_inst_dmem_n1770,
         mem_stage_inst_dmem_n1769, mem_stage_inst_dmem_n1768,
         mem_stage_inst_dmem_n1767, mem_stage_inst_dmem_n1766,
         mem_stage_inst_dmem_n1765, mem_stage_inst_dmem_n1764,
         mem_stage_inst_dmem_n1763, mem_stage_inst_dmem_n1762,
         mem_stage_inst_dmem_n1761, mem_stage_inst_dmem_n1760,
         mem_stage_inst_dmem_n1759, mem_stage_inst_dmem_n1758,
         mem_stage_inst_dmem_n1757, mem_stage_inst_dmem_n1756,
         mem_stage_inst_dmem_n1755, mem_stage_inst_dmem_n1754,
         mem_stage_inst_dmem_n1753, mem_stage_inst_dmem_n1752,
         mem_stage_inst_dmem_n1751, mem_stage_inst_dmem_n1750,
         mem_stage_inst_dmem_n1749, mem_stage_inst_dmem_n1748,
         mem_stage_inst_dmem_n1747, mem_stage_inst_dmem_n1746,
         mem_stage_inst_dmem_n1745, mem_stage_inst_dmem_n1744,
         mem_stage_inst_dmem_n1743, mem_stage_inst_dmem_n1742,
         mem_stage_inst_dmem_n1741, mem_stage_inst_dmem_n1740,
         mem_stage_inst_dmem_n1739, mem_stage_inst_dmem_n1738,
         mem_stage_inst_dmem_n1737, mem_stage_inst_dmem_n1736,
         mem_stage_inst_dmem_n1735, mem_stage_inst_dmem_n1734,
         mem_stage_inst_dmem_n1733, mem_stage_inst_dmem_n1732,
         mem_stage_inst_dmem_n1731, mem_stage_inst_dmem_n1730,
         mem_stage_inst_dmem_n1729, mem_stage_inst_dmem_n1728,
         mem_stage_inst_dmem_n1727, mem_stage_inst_dmem_n1726,
         mem_stage_inst_dmem_n1725, mem_stage_inst_dmem_n1724,
         mem_stage_inst_dmem_n1723, mem_stage_inst_dmem_n1722,
         mem_stage_inst_dmem_n1721, mem_stage_inst_dmem_n1720,
         mem_stage_inst_dmem_n1719, mem_stage_inst_dmem_n1718,
         mem_stage_inst_dmem_n1717, mem_stage_inst_dmem_n1716,
         mem_stage_inst_dmem_n1715, mem_stage_inst_dmem_n1714,
         mem_stage_inst_dmem_n1713, mem_stage_inst_dmem_n1712,
         mem_stage_inst_dmem_n1711, mem_stage_inst_dmem_n1710,
         mem_stage_inst_dmem_n1709, mem_stage_inst_dmem_n1708,
         mem_stage_inst_dmem_n1707, mem_stage_inst_dmem_n1706,
         mem_stage_inst_dmem_n1705, mem_stage_inst_dmem_n1704,
         mem_stage_inst_dmem_n1703, mem_stage_inst_dmem_n1702,
         mem_stage_inst_dmem_n1701, mem_stage_inst_dmem_n1700,
         mem_stage_inst_dmem_n1699, mem_stage_inst_dmem_n1698,
         mem_stage_inst_dmem_n1697, mem_stage_inst_dmem_n1696,
         mem_stage_inst_dmem_n1695, mem_stage_inst_dmem_n1694,
         mem_stage_inst_dmem_n1693, mem_stage_inst_dmem_n1692,
         mem_stage_inst_dmem_n1691, mem_stage_inst_dmem_n1690,
         mem_stage_inst_dmem_n1689, mem_stage_inst_dmem_n1688,
         mem_stage_inst_dmem_n1687, mem_stage_inst_dmem_n1686,
         mem_stage_inst_dmem_n1685, mem_stage_inst_dmem_n1684,
         mem_stage_inst_dmem_n1683, mem_stage_inst_dmem_n1682,
         mem_stage_inst_dmem_n1681, mem_stage_inst_dmem_n1680,
         mem_stage_inst_dmem_n1679, mem_stage_inst_dmem_n1678,
         mem_stage_inst_dmem_n1677, mem_stage_inst_dmem_n1676,
         mem_stage_inst_dmem_n1675, mem_stage_inst_dmem_n1674,
         mem_stage_inst_dmem_n1673, mem_stage_inst_dmem_n1672,
         mem_stage_inst_dmem_n1671, mem_stage_inst_dmem_n1670,
         mem_stage_inst_dmem_n1669, mem_stage_inst_dmem_n1668,
         mem_stage_inst_dmem_n1667, mem_stage_inst_dmem_n1666,
         mem_stage_inst_dmem_n1665, mem_stage_inst_dmem_n1664,
         mem_stage_inst_dmem_n1663, mem_stage_inst_dmem_n1662,
         mem_stage_inst_dmem_n1661, mem_stage_inst_dmem_n1660,
         mem_stage_inst_dmem_n1659, mem_stage_inst_dmem_n1658,
         mem_stage_inst_dmem_n1657, mem_stage_inst_dmem_n1656,
         mem_stage_inst_dmem_n1655, mem_stage_inst_dmem_n1654,
         mem_stage_inst_dmem_n1653, mem_stage_inst_dmem_n1652,
         mem_stage_inst_dmem_n1651, mem_stage_inst_dmem_n1650,
         mem_stage_inst_dmem_n1649, mem_stage_inst_dmem_n1648,
         mem_stage_inst_dmem_n1647, mem_stage_inst_dmem_n1646,
         mem_stage_inst_dmem_n1645, mem_stage_inst_dmem_n1644,
         mem_stage_inst_dmem_n1643, mem_stage_inst_dmem_n1642,
         mem_stage_inst_dmem_n1641, mem_stage_inst_dmem_n1640,
         mem_stage_inst_dmem_n1639, mem_stage_inst_dmem_n1638,
         mem_stage_inst_dmem_n1637, mem_stage_inst_dmem_n1636,
         mem_stage_inst_dmem_n1635, mem_stage_inst_dmem_n1634,
         mem_stage_inst_dmem_n1633, mem_stage_inst_dmem_n1632,
         mem_stage_inst_dmem_n1631, mem_stage_inst_dmem_n1630,
         mem_stage_inst_dmem_n1629, mem_stage_inst_dmem_n1628,
         mem_stage_inst_dmem_n1627, mem_stage_inst_dmem_n1626,
         mem_stage_inst_dmem_n1625, mem_stage_inst_dmem_n1624,
         mem_stage_inst_dmem_n1623, mem_stage_inst_dmem_n1622,
         mem_stage_inst_dmem_n1621, mem_stage_inst_dmem_n1620,
         mem_stage_inst_dmem_n1619, mem_stage_inst_dmem_n1618,
         mem_stage_inst_dmem_n1617, mem_stage_inst_dmem_n1616,
         mem_stage_inst_dmem_n1615, mem_stage_inst_dmem_n1614,
         mem_stage_inst_dmem_n1613, mem_stage_inst_dmem_n1612,
         mem_stage_inst_dmem_n1611, mem_stage_inst_dmem_n1610,
         mem_stage_inst_dmem_n1609, mem_stage_inst_dmem_n1608,
         mem_stage_inst_dmem_n1607, mem_stage_inst_dmem_n1606,
         mem_stage_inst_dmem_n1605, mem_stage_inst_dmem_n1604,
         mem_stage_inst_dmem_n1603, mem_stage_inst_dmem_n1602,
         mem_stage_inst_dmem_n1601, mem_stage_inst_dmem_n1600,
         mem_stage_inst_dmem_n1599, mem_stage_inst_dmem_n1598,
         mem_stage_inst_dmem_n1597, mem_stage_inst_dmem_n1596,
         mem_stage_inst_dmem_n1595, mem_stage_inst_dmem_n1594,
         mem_stage_inst_dmem_n1593, mem_stage_inst_dmem_n1592,
         mem_stage_inst_dmem_n1591, mem_stage_inst_dmem_n1590,
         mem_stage_inst_dmem_n1589, mem_stage_inst_dmem_n1588,
         mem_stage_inst_dmem_n1587, mem_stage_inst_dmem_n1586,
         mem_stage_inst_dmem_n1585, mem_stage_inst_dmem_n1584,
         mem_stage_inst_dmem_n1583, mem_stage_inst_dmem_n1582,
         mem_stage_inst_dmem_n1581, mem_stage_inst_dmem_n1580,
         mem_stage_inst_dmem_n1579, mem_stage_inst_dmem_n1578,
         mem_stage_inst_dmem_n1577, mem_stage_inst_dmem_n1576,
         mem_stage_inst_dmem_n1575, mem_stage_inst_dmem_n1574,
         mem_stage_inst_dmem_n1573, mem_stage_inst_dmem_n1572,
         mem_stage_inst_dmem_n1571, mem_stage_inst_dmem_n1570,
         mem_stage_inst_dmem_n1569, mem_stage_inst_dmem_n1568,
         mem_stage_inst_dmem_n1567, mem_stage_inst_dmem_n1566,
         mem_stage_inst_dmem_n1565, mem_stage_inst_dmem_n1564,
         mem_stage_inst_dmem_n1563, mem_stage_inst_dmem_n1562,
         mem_stage_inst_dmem_n1561, mem_stage_inst_dmem_n1560,
         mem_stage_inst_dmem_n1559, mem_stage_inst_dmem_n1558,
         mem_stage_inst_dmem_n1557, mem_stage_inst_dmem_n1556,
         mem_stage_inst_dmem_n1555, mem_stage_inst_dmem_n1554,
         mem_stage_inst_dmem_n1553, mem_stage_inst_dmem_n1552,
         mem_stage_inst_dmem_n1551, mem_stage_inst_dmem_n1550,
         mem_stage_inst_dmem_n1549, mem_stage_inst_dmem_n1548,
         mem_stage_inst_dmem_n1547, mem_stage_inst_dmem_n1546,
         mem_stage_inst_dmem_n1545, mem_stage_inst_dmem_n1544,
         mem_stage_inst_dmem_n1543, mem_stage_inst_dmem_n1542,
         mem_stage_inst_dmem_n1541, mem_stage_inst_dmem_n1540,
         mem_stage_inst_dmem_n1539, mem_stage_inst_dmem_n1538,
         mem_stage_inst_dmem_n1537, mem_stage_inst_dmem_n1536,
         mem_stage_inst_dmem_n1535, mem_stage_inst_dmem_n1534,
         mem_stage_inst_dmem_n1533, mem_stage_inst_dmem_n1532,
         mem_stage_inst_dmem_n1531, mem_stage_inst_dmem_n1530,
         mem_stage_inst_dmem_n1529, mem_stage_inst_dmem_n1528,
         mem_stage_inst_dmem_n1527, mem_stage_inst_dmem_n1526,
         mem_stage_inst_dmem_n1525, mem_stage_inst_dmem_n1524,
         mem_stage_inst_dmem_n1523, mem_stage_inst_dmem_n1522,
         mem_stage_inst_dmem_n1521, mem_stage_inst_dmem_n1520,
         mem_stage_inst_dmem_n1519, mem_stage_inst_dmem_n1518,
         mem_stage_inst_dmem_n1517, mem_stage_inst_dmem_n1516,
         mem_stage_inst_dmem_n1515, mem_stage_inst_dmem_n1514,
         mem_stage_inst_dmem_n1513, mem_stage_inst_dmem_n1512,
         mem_stage_inst_dmem_n1511, mem_stage_inst_dmem_n1510,
         mem_stage_inst_dmem_n1509, mem_stage_inst_dmem_n1508,
         mem_stage_inst_dmem_n1507, mem_stage_inst_dmem_n1506,
         mem_stage_inst_dmem_n1505, mem_stage_inst_dmem_n1504,
         mem_stage_inst_dmem_n1503, mem_stage_inst_dmem_n1502,
         mem_stage_inst_dmem_n1501, mem_stage_inst_dmem_n1500,
         mem_stage_inst_dmem_n1499, mem_stage_inst_dmem_n1498,
         mem_stage_inst_dmem_n1497, mem_stage_inst_dmem_n1496,
         mem_stage_inst_dmem_n1495, mem_stage_inst_dmem_n1494,
         mem_stage_inst_dmem_n1493, mem_stage_inst_dmem_n1492,
         mem_stage_inst_dmem_n1491, mem_stage_inst_dmem_n1490,
         mem_stage_inst_dmem_n1489, mem_stage_inst_dmem_n1488,
         mem_stage_inst_dmem_n1487, mem_stage_inst_dmem_n1486,
         mem_stage_inst_dmem_n1485, mem_stage_inst_dmem_n1484,
         mem_stage_inst_dmem_n1483, mem_stage_inst_dmem_n1482,
         mem_stage_inst_dmem_n1481, mem_stage_inst_dmem_n1480,
         mem_stage_inst_dmem_n1479, mem_stage_inst_dmem_n1478,
         mem_stage_inst_dmem_n1477, mem_stage_inst_dmem_n1476,
         mem_stage_inst_dmem_n1475, mem_stage_inst_dmem_n1474,
         mem_stage_inst_dmem_n1473, mem_stage_inst_dmem_n1472,
         mem_stage_inst_dmem_n1471, mem_stage_inst_dmem_n1470,
         mem_stage_inst_dmem_n1469, mem_stage_inst_dmem_n1468,
         mem_stage_inst_dmem_n1467, mem_stage_inst_dmem_n1466,
         mem_stage_inst_dmem_n1465, mem_stage_inst_dmem_n1464,
         mem_stage_inst_dmem_n1463, mem_stage_inst_dmem_n1462,
         mem_stage_inst_dmem_n1461, mem_stage_inst_dmem_n1460,
         mem_stage_inst_dmem_n1459, mem_stage_inst_dmem_n1458,
         mem_stage_inst_dmem_n1457, mem_stage_inst_dmem_n1456,
         mem_stage_inst_dmem_n1455, mem_stage_inst_dmem_n1454,
         mem_stage_inst_dmem_n1453, mem_stage_inst_dmem_n1452,
         mem_stage_inst_dmem_n1451, mem_stage_inst_dmem_n1450,
         mem_stage_inst_dmem_n1449, mem_stage_inst_dmem_n1448,
         mem_stage_inst_dmem_n1447, mem_stage_inst_dmem_n1446,
         mem_stage_inst_dmem_n1445, mem_stage_inst_dmem_n1444,
         mem_stage_inst_dmem_n1443, mem_stage_inst_dmem_n1442,
         mem_stage_inst_dmem_n1441, mem_stage_inst_dmem_n1440,
         mem_stage_inst_dmem_n1439, mem_stage_inst_dmem_n1438,
         mem_stage_inst_dmem_n1437, mem_stage_inst_dmem_n1436,
         mem_stage_inst_dmem_n1435, mem_stage_inst_dmem_n1434,
         mem_stage_inst_dmem_n1433, mem_stage_inst_dmem_n1432,
         mem_stage_inst_dmem_n1431, mem_stage_inst_dmem_n1430,
         mem_stage_inst_dmem_n1429, mem_stage_inst_dmem_n1428,
         mem_stage_inst_dmem_n1427, mem_stage_inst_dmem_n1426,
         mem_stage_inst_dmem_n1425, mem_stage_inst_dmem_n1424,
         mem_stage_inst_dmem_n1423, mem_stage_inst_dmem_n1422,
         mem_stage_inst_dmem_n1421, mem_stage_inst_dmem_n1420,
         mem_stage_inst_dmem_n1419, mem_stage_inst_dmem_n1418,
         mem_stage_inst_dmem_n1417, mem_stage_inst_dmem_n1416,
         mem_stage_inst_dmem_n1415, mem_stage_inst_dmem_n1414,
         mem_stage_inst_dmem_n1413, mem_stage_inst_dmem_n1412,
         mem_stage_inst_dmem_n1411, mem_stage_inst_dmem_n1410,
         mem_stage_inst_dmem_n1409, mem_stage_inst_dmem_n1408,
         mem_stage_inst_dmem_n1407, mem_stage_inst_dmem_n1406,
         mem_stage_inst_dmem_n1405, mem_stage_inst_dmem_n1404,
         mem_stage_inst_dmem_n1403, mem_stage_inst_dmem_n1402,
         mem_stage_inst_dmem_n1401, mem_stage_inst_dmem_n1400,
         mem_stage_inst_dmem_n1399, mem_stage_inst_dmem_n1398,
         mem_stage_inst_dmem_n1397, mem_stage_inst_dmem_n1396,
         mem_stage_inst_dmem_n1395, mem_stage_inst_dmem_n1394,
         mem_stage_inst_dmem_n1393, mem_stage_inst_dmem_n1392,
         mem_stage_inst_dmem_n1391, mem_stage_inst_dmem_n1390,
         mem_stage_inst_dmem_n1389, mem_stage_inst_dmem_n1388,
         mem_stage_inst_dmem_n1387, mem_stage_inst_dmem_n1386,
         mem_stage_inst_dmem_n1385, mem_stage_inst_dmem_n1384,
         mem_stage_inst_dmem_n1383, mem_stage_inst_dmem_n1382,
         mem_stage_inst_dmem_n1381, mem_stage_inst_dmem_n1380,
         mem_stage_inst_dmem_n1379, mem_stage_inst_dmem_n1378,
         mem_stage_inst_dmem_n1377, mem_stage_inst_dmem_n1376,
         mem_stage_inst_dmem_n1375, mem_stage_inst_dmem_n1374,
         mem_stage_inst_dmem_n1373, mem_stage_inst_dmem_n1372,
         mem_stage_inst_dmem_n1371, mem_stage_inst_dmem_n1370,
         mem_stage_inst_dmem_n1369, mem_stage_inst_dmem_n1368,
         mem_stage_inst_dmem_n1367, mem_stage_inst_dmem_n1366,
         mem_stage_inst_dmem_n1365, mem_stage_inst_dmem_n1364,
         mem_stage_inst_dmem_n1363, mem_stage_inst_dmem_n1362,
         mem_stage_inst_dmem_n1361, mem_stage_inst_dmem_n1360,
         mem_stage_inst_dmem_n1359, mem_stage_inst_dmem_n1358,
         mem_stage_inst_dmem_n1357, mem_stage_inst_dmem_n1356,
         mem_stage_inst_dmem_n1355, mem_stage_inst_dmem_n1354,
         mem_stage_inst_dmem_n1353, mem_stage_inst_dmem_n1352,
         mem_stage_inst_dmem_n1351, mem_stage_inst_dmem_n1350,
         mem_stage_inst_dmem_n1349, mem_stage_inst_dmem_n1348,
         mem_stage_inst_dmem_n1347, mem_stage_inst_dmem_n1346,
         mem_stage_inst_dmem_n1345, mem_stage_inst_dmem_n1344,
         mem_stage_inst_dmem_n1343, mem_stage_inst_dmem_n1342,
         mem_stage_inst_dmem_n1341, mem_stage_inst_dmem_n1340,
         mem_stage_inst_dmem_n1339, mem_stage_inst_dmem_n1338,
         mem_stage_inst_dmem_n1337, mem_stage_inst_dmem_n1336,
         mem_stage_inst_dmem_n1335, mem_stage_inst_dmem_n1334,
         mem_stage_inst_dmem_n1333, mem_stage_inst_dmem_n1332,
         mem_stage_inst_dmem_n1331, mem_stage_inst_dmem_n1330,
         mem_stage_inst_dmem_n1329, mem_stage_inst_dmem_n1328,
         mem_stage_inst_dmem_n1327, mem_stage_inst_dmem_n1326,
         mem_stage_inst_dmem_n1325, mem_stage_inst_dmem_n1324,
         mem_stage_inst_dmem_n1323, mem_stage_inst_dmem_n1322,
         mem_stage_inst_dmem_n1321, mem_stage_inst_dmem_n1320,
         mem_stage_inst_dmem_n1319, mem_stage_inst_dmem_n1318,
         mem_stage_inst_dmem_n1317, mem_stage_inst_dmem_n1316,
         mem_stage_inst_dmem_n1315, mem_stage_inst_dmem_n1314,
         mem_stage_inst_dmem_n1313, mem_stage_inst_dmem_n1312,
         mem_stage_inst_dmem_n1311, mem_stage_inst_dmem_n1310,
         mem_stage_inst_dmem_n1309, mem_stage_inst_dmem_n1308,
         mem_stage_inst_dmem_n1307, mem_stage_inst_dmem_n1306,
         mem_stage_inst_dmem_n1305, mem_stage_inst_dmem_n1304,
         mem_stage_inst_dmem_n1303, mem_stage_inst_dmem_n1302,
         mem_stage_inst_dmem_n1301, mem_stage_inst_dmem_n1300,
         mem_stage_inst_dmem_n1299, mem_stage_inst_dmem_n1298,
         mem_stage_inst_dmem_n1297, mem_stage_inst_dmem_n1296,
         mem_stage_inst_dmem_n1295, mem_stage_inst_dmem_n1294,
         mem_stage_inst_dmem_n1293, mem_stage_inst_dmem_n1292,
         mem_stage_inst_dmem_n1291, mem_stage_inst_dmem_n1290,
         mem_stage_inst_dmem_n1289, mem_stage_inst_dmem_n1288,
         mem_stage_inst_dmem_n1287, mem_stage_inst_dmem_n1286,
         mem_stage_inst_dmem_n1285, mem_stage_inst_dmem_n1284,
         mem_stage_inst_dmem_n1283, mem_stage_inst_dmem_n1282,
         mem_stage_inst_dmem_n1281, mem_stage_inst_dmem_n1280,
         mem_stage_inst_dmem_n1279, mem_stage_inst_dmem_n1278,
         mem_stage_inst_dmem_n1277, mem_stage_inst_dmem_n1276,
         mem_stage_inst_dmem_n1275, mem_stage_inst_dmem_n1274,
         mem_stage_inst_dmem_n1273, mem_stage_inst_dmem_n1272,
         mem_stage_inst_dmem_n1271, mem_stage_inst_dmem_n1270,
         mem_stage_inst_dmem_n1269, mem_stage_inst_dmem_n1268,
         mem_stage_inst_dmem_n1267, mem_stage_inst_dmem_n1266,
         mem_stage_inst_dmem_n1265, mem_stage_inst_dmem_n1264,
         mem_stage_inst_dmem_n1263, mem_stage_inst_dmem_n1262,
         mem_stage_inst_dmem_n1261, mem_stage_inst_dmem_n1260,
         mem_stage_inst_dmem_n1259, mem_stage_inst_dmem_n1258,
         mem_stage_inst_dmem_n1257, mem_stage_inst_dmem_n1256,
         mem_stage_inst_dmem_n1255, mem_stage_inst_dmem_n1254,
         mem_stage_inst_dmem_n1253, mem_stage_inst_dmem_n1252,
         mem_stage_inst_dmem_n1251, mem_stage_inst_dmem_n1250,
         mem_stage_inst_dmem_n1249, mem_stage_inst_dmem_n1248,
         mem_stage_inst_dmem_n1247, mem_stage_inst_dmem_n1246,
         mem_stage_inst_dmem_n1245, mem_stage_inst_dmem_n1244,
         mem_stage_inst_dmem_n1243, mem_stage_inst_dmem_n1242,
         mem_stage_inst_dmem_n1241, mem_stage_inst_dmem_n1240,
         mem_stage_inst_dmem_n1239, mem_stage_inst_dmem_n1238,
         mem_stage_inst_dmem_n1237, mem_stage_inst_dmem_n1236,
         mem_stage_inst_dmem_n1235, mem_stage_inst_dmem_n1234,
         mem_stage_inst_dmem_n1233, mem_stage_inst_dmem_n1232,
         mem_stage_inst_dmem_n1231, mem_stage_inst_dmem_n1230,
         mem_stage_inst_dmem_n1229, mem_stage_inst_dmem_n1228,
         mem_stage_inst_dmem_n1227, mem_stage_inst_dmem_n1226,
         mem_stage_inst_dmem_n1225, mem_stage_inst_dmem_n1224,
         mem_stage_inst_dmem_n1223, mem_stage_inst_dmem_n1222,
         mem_stage_inst_dmem_n1221, mem_stage_inst_dmem_n1220,
         mem_stage_inst_dmem_n1219, mem_stage_inst_dmem_n1218,
         mem_stage_inst_dmem_n1217, mem_stage_inst_dmem_n1216,
         mem_stage_inst_dmem_n1215, mem_stage_inst_dmem_n1214,
         mem_stage_inst_dmem_n1213, mem_stage_inst_dmem_n1212,
         mem_stage_inst_dmem_n1211, mem_stage_inst_dmem_n1210,
         mem_stage_inst_dmem_n1209, mem_stage_inst_dmem_n1208,
         mem_stage_inst_dmem_n1207, mem_stage_inst_dmem_n1206,
         mem_stage_inst_dmem_n1205, mem_stage_inst_dmem_n1204,
         mem_stage_inst_dmem_n1203, mem_stage_inst_dmem_n1202,
         mem_stage_inst_dmem_n1201, mem_stage_inst_dmem_n1200,
         mem_stage_inst_dmem_n1199, mem_stage_inst_dmem_n1198,
         mem_stage_inst_dmem_n1197, mem_stage_inst_dmem_n1196,
         mem_stage_inst_dmem_n1195, mem_stage_inst_dmem_n1194,
         mem_stage_inst_dmem_n1193, mem_stage_inst_dmem_n1192,
         mem_stage_inst_dmem_n1191, mem_stage_inst_dmem_n1190,
         mem_stage_inst_dmem_n1189, mem_stage_inst_dmem_n1188,
         mem_stage_inst_dmem_n1187, mem_stage_inst_dmem_n1186,
         mem_stage_inst_dmem_n1185, mem_stage_inst_dmem_n1184,
         mem_stage_inst_dmem_n1183, mem_stage_inst_dmem_n1182,
         mem_stage_inst_dmem_n1181, mem_stage_inst_dmem_n1180,
         mem_stage_inst_dmem_n1179, mem_stage_inst_dmem_n1178,
         mem_stage_inst_dmem_n1177, mem_stage_inst_dmem_n1176,
         mem_stage_inst_dmem_n1175, mem_stage_inst_dmem_n1174,
         mem_stage_inst_dmem_n1173, mem_stage_inst_dmem_n1172,
         mem_stage_inst_dmem_n1171, mem_stage_inst_dmem_n1170,
         mem_stage_inst_dmem_n1169, mem_stage_inst_dmem_n1168,
         mem_stage_inst_dmem_n1167, mem_stage_inst_dmem_n1166,
         mem_stage_inst_dmem_n1165, mem_stage_inst_dmem_n1164,
         mem_stage_inst_dmem_n1163, mem_stage_inst_dmem_n1162,
         mem_stage_inst_dmem_n1161, mem_stage_inst_dmem_n1160,
         mem_stage_inst_dmem_n1159, mem_stage_inst_dmem_n1158,
         mem_stage_inst_dmem_n1157, mem_stage_inst_dmem_n1156,
         mem_stage_inst_dmem_n1155, mem_stage_inst_dmem_n1154,
         mem_stage_inst_dmem_n1153, mem_stage_inst_dmem_n1152,
         mem_stage_inst_dmem_n1151, mem_stage_inst_dmem_n1150,
         mem_stage_inst_dmem_n1149, mem_stage_inst_dmem_n1148,
         mem_stage_inst_dmem_n1147, mem_stage_inst_dmem_n1146,
         mem_stage_inst_dmem_n1145, mem_stage_inst_dmem_n1144,
         mem_stage_inst_dmem_n1143, mem_stage_inst_dmem_n1142,
         mem_stage_inst_dmem_n1141, mem_stage_inst_dmem_n1140,
         mem_stage_inst_dmem_n1139, mem_stage_inst_dmem_n1138,
         mem_stage_inst_dmem_n1137, mem_stage_inst_dmem_n1136,
         mem_stage_inst_dmem_n1135, mem_stage_inst_dmem_n1134,
         mem_stage_inst_dmem_n1133, mem_stage_inst_dmem_n1132,
         mem_stage_inst_dmem_n1131, mem_stage_inst_dmem_n1130,
         mem_stage_inst_dmem_n1129, mem_stage_inst_dmem_n1128,
         mem_stage_inst_dmem_n1127, mem_stage_inst_dmem_n1126,
         mem_stage_inst_dmem_n1125, mem_stage_inst_dmem_n1124,
         mem_stage_inst_dmem_n1123, mem_stage_inst_dmem_n1122,
         mem_stage_inst_dmem_n1121, mem_stage_inst_dmem_n1120,
         mem_stage_inst_dmem_n1119, mem_stage_inst_dmem_n1118,
         mem_stage_inst_dmem_n1117, mem_stage_inst_dmem_n1116,
         mem_stage_inst_dmem_n1115, mem_stage_inst_dmem_n1114,
         mem_stage_inst_dmem_n1113, mem_stage_inst_dmem_n1112,
         mem_stage_inst_dmem_n1111, mem_stage_inst_dmem_n1110,
         mem_stage_inst_dmem_n1109, mem_stage_inst_dmem_n1108,
         mem_stage_inst_dmem_n1107, mem_stage_inst_dmem_n1106,
         mem_stage_inst_dmem_n1105, mem_stage_inst_dmem_n1104,
         mem_stage_inst_dmem_n1103, mem_stage_inst_dmem_n1102,
         mem_stage_inst_dmem_n1101, mem_stage_inst_dmem_n1100,
         mem_stage_inst_dmem_n1099, mem_stage_inst_dmem_n1098,
         mem_stage_inst_dmem_n1097, mem_stage_inst_dmem_n1096,
         mem_stage_inst_dmem_n1095, mem_stage_inst_dmem_n1094,
         mem_stage_inst_dmem_n1093, mem_stage_inst_dmem_n1092,
         mem_stage_inst_dmem_n1091, mem_stage_inst_dmem_n1090,
         mem_stage_inst_dmem_n1089, mem_stage_inst_dmem_n1088,
         mem_stage_inst_dmem_n1087, mem_stage_inst_dmem_n1086,
         mem_stage_inst_dmem_n1085, mem_stage_inst_dmem_n1084,
         mem_stage_inst_dmem_n1083, mem_stage_inst_dmem_n1082,
         mem_stage_inst_dmem_n1081, mem_stage_inst_dmem_n1080,
         mem_stage_inst_dmem_n1079, mem_stage_inst_dmem_n1078,
         mem_stage_inst_dmem_n1077, mem_stage_inst_dmem_n1076,
         mem_stage_inst_dmem_n1075, mem_stage_inst_dmem_n1074,
         mem_stage_inst_dmem_n1073, mem_stage_inst_dmem_n1072,
         mem_stage_inst_dmem_n1071, mem_stage_inst_dmem_n1070,
         mem_stage_inst_dmem_n1069, mem_stage_inst_dmem_n1068,
         mem_stage_inst_dmem_n1067, mem_stage_inst_dmem_n1066,
         mem_stage_inst_dmem_n1065, mem_stage_inst_dmem_n1064,
         mem_stage_inst_dmem_n1063, mem_stage_inst_dmem_n1062,
         mem_stage_inst_dmem_n1061, mem_stage_inst_dmem_n1060,
         mem_stage_inst_dmem_n1059, mem_stage_inst_dmem_n1058,
         mem_stage_inst_dmem_n1057, mem_stage_inst_dmem_n1056,
         mem_stage_inst_dmem_n1055, mem_stage_inst_dmem_n1054,
         mem_stage_inst_dmem_n1053, mem_stage_inst_dmem_n1052,
         mem_stage_inst_dmem_n1051, mem_stage_inst_dmem_n1050,
         mem_stage_inst_dmem_n1049, mem_stage_inst_dmem_n1048,
         mem_stage_inst_dmem_n1047, mem_stage_inst_dmem_n1046,
         mem_stage_inst_dmem_n1045, mem_stage_inst_dmem_n1044,
         mem_stage_inst_dmem_n1043, mem_stage_inst_dmem_n1042,
         mem_stage_inst_dmem_n1041, mem_stage_inst_dmem_n1040,
         mem_stage_inst_dmem_n1039, mem_stage_inst_dmem_n1038,
         mem_stage_inst_dmem_n1037, mem_stage_inst_dmem_n1036,
         mem_stage_inst_dmem_n1035, mem_stage_inst_dmem_n1034,
         mem_stage_inst_dmem_n1033, mem_stage_inst_dmem_n1032,
         mem_stage_inst_dmem_n1031, mem_stage_inst_dmem_n1030,
         mem_stage_inst_dmem_n1029, mem_stage_inst_dmem_n1028,
         mem_stage_inst_dmem_n1027, mem_stage_inst_dmem_n1026,
         mem_stage_inst_dmem_n1025, mem_stage_inst_dmem_n1024,
         mem_stage_inst_dmem_n1023, mem_stage_inst_dmem_n1022,
         mem_stage_inst_dmem_n1021, mem_stage_inst_dmem_n1020,
         mem_stage_inst_dmem_n1019, mem_stage_inst_dmem_n1018,
         mem_stage_inst_dmem_n1017, mem_stage_inst_dmem_n1016,
         mem_stage_inst_dmem_n1015, mem_stage_inst_dmem_n1014,
         mem_stage_inst_dmem_n1013, mem_stage_inst_dmem_n1012,
         mem_stage_inst_dmem_n1011, mem_stage_inst_dmem_n1010,
         mem_stage_inst_dmem_n1009, mem_stage_inst_dmem_n1008,
         mem_stage_inst_dmem_n1007, mem_stage_inst_dmem_n1006,
         mem_stage_inst_dmem_n1005, mem_stage_inst_dmem_n1004,
         mem_stage_inst_dmem_n1003, mem_stage_inst_dmem_n1002,
         mem_stage_inst_dmem_n1001, mem_stage_inst_dmem_n1000,
         mem_stage_inst_dmem_n999, mem_stage_inst_dmem_n998,
         mem_stage_inst_dmem_n997, mem_stage_inst_dmem_n996,
         mem_stage_inst_dmem_n995, mem_stage_inst_dmem_n994,
         mem_stage_inst_dmem_n993, mem_stage_inst_dmem_n992,
         mem_stage_inst_dmem_n991, mem_stage_inst_dmem_n990,
         mem_stage_inst_dmem_n989, mem_stage_inst_dmem_n988,
         mem_stage_inst_dmem_n987, mem_stage_inst_dmem_n986,
         mem_stage_inst_dmem_n985, mem_stage_inst_dmem_n984,
         mem_stage_inst_dmem_n983, mem_stage_inst_dmem_n982,
         mem_stage_inst_dmem_n981, mem_stage_inst_dmem_n980,
         mem_stage_inst_dmem_n979, mem_stage_inst_dmem_n978,
         mem_stage_inst_dmem_n977, mem_stage_inst_dmem_n976,
         mem_stage_inst_dmem_n975, mem_stage_inst_dmem_n974,
         mem_stage_inst_dmem_n973, mem_stage_inst_dmem_n972,
         mem_stage_inst_dmem_n971, mem_stage_inst_dmem_n970,
         mem_stage_inst_dmem_n969, mem_stage_inst_dmem_n968,
         mem_stage_inst_dmem_n967, mem_stage_inst_dmem_n966,
         mem_stage_inst_dmem_n965, mem_stage_inst_dmem_n964,
         mem_stage_inst_dmem_n963, mem_stage_inst_dmem_n962,
         mem_stage_inst_dmem_n961, mem_stage_inst_dmem_n960,
         mem_stage_inst_dmem_n959, mem_stage_inst_dmem_n958,
         mem_stage_inst_dmem_n957, mem_stage_inst_dmem_n956,
         mem_stage_inst_dmem_n955, mem_stage_inst_dmem_n954,
         mem_stage_inst_dmem_n953, mem_stage_inst_dmem_n952,
         mem_stage_inst_dmem_n951, mem_stage_inst_dmem_n950,
         mem_stage_inst_dmem_n949, mem_stage_inst_dmem_n948,
         mem_stage_inst_dmem_n947, mem_stage_inst_dmem_n946,
         mem_stage_inst_dmem_n945, mem_stage_inst_dmem_n944,
         mem_stage_inst_dmem_n943, mem_stage_inst_dmem_n942,
         mem_stage_inst_dmem_n941, mem_stage_inst_dmem_n940,
         mem_stage_inst_dmem_n939, mem_stage_inst_dmem_n938,
         mem_stage_inst_dmem_n937, mem_stage_inst_dmem_n936,
         mem_stage_inst_dmem_n935, mem_stage_inst_dmem_n934,
         mem_stage_inst_dmem_n933, mem_stage_inst_dmem_n932,
         mem_stage_inst_dmem_n931, mem_stage_inst_dmem_n930,
         mem_stage_inst_dmem_n929, mem_stage_inst_dmem_n928,
         mem_stage_inst_dmem_n927, mem_stage_inst_dmem_n926,
         mem_stage_inst_dmem_n925, mem_stage_inst_dmem_n924,
         mem_stage_inst_dmem_n923, mem_stage_inst_dmem_n922,
         mem_stage_inst_dmem_n921, mem_stage_inst_dmem_n920,
         mem_stage_inst_dmem_n919, mem_stage_inst_dmem_n918,
         mem_stage_inst_dmem_n917, mem_stage_inst_dmem_n916,
         mem_stage_inst_dmem_n915, mem_stage_inst_dmem_n914,
         mem_stage_inst_dmem_n913, mem_stage_inst_dmem_n912,
         mem_stage_inst_dmem_n911, mem_stage_inst_dmem_n910,
         mem_stage_inst_dmem_n909, mem_stage_inst_dmem_n908,
         mem_stage_inst_dmem_n907, mem_stage_inst_dmem_n906,
         mem_stage_inst_dmem_n905, mem_stage_inst_dmem_n904,
         mem_stage_inst_dmem_n903, mem_stage_inst_dmem_n902,
         mem_stage_inst_dmem_n901, mem_stage_inst_dmem_n900,
         mem_stage_inst_dmem_n899, mem_stage_inst_dmem_n898,
         mem_stage_inst_dmem_n897, mem_stage_inst_dmem_n896,
         mem_stage_inst_dmem_n895, mem_stage_inst_dmem_n894,
         mem_stage_inst_dmem_n893, mem_stage_inst_dmem_n892,
         mem_stage_inst_dmem_n891, mem_stage_inst_dmem_n890,
         mem_stage_inst_dmem_n889, mem_stage_inst_dmem_n888,
         mem_stage_inst_dmem_n887, mem_stage_inst_dmem_n886,
         mem_stage_inst_dmem_n885, mem_stage_inst_dmem_n884,
         mem_stage_inst_dmem_n883, mem_stage_inst_dmem_n882,
         mem_stage_inst_dmem_n881, mem_stage_inst_dmem_n880,
         mem_stage_inst_dmem_n879, mem_stage_inst_dmem_n878,
         mem_stage_inst_dmem_n877, mem_stage_inst_dmem_n876,
         mem_stage_inst_dmem_n875, mem_stage_inst_dmem_n874,
         mem_stage_inst_dmem_n873, mem_stage_inst_dmem_n872,
         mem_stage_inst_dmem_n871, mem_stage_inst_dmem_n870,
         mem_stage_inst_dmem_n869, mem_stage_inst_dmem_n868,
         mem_stage_inst_dmem_n867, mem_stage_inst_dmem_n866,
         mem_stage_inst_dmem_n865, mem_stage_inst_dmem_n864,
         mem_stage_inst_dmem_n863, mem_stage_inst_dmem_n862,
         mem_stage_inst_dmem_n861, mem_stage_inst_dmem_n860,
         mem_stage_inst_dmem_n859, mem_stage_inst_dmem_n858,
         mem_stage_inst_dmem_n857, mem_stage_inst_dmem_n856,
         mem_stage_inst_dmem_n855, mem_stage_inst_dmem_n854,
         mem_stage_inst_dmem_n853, mem_stage_inst_dmem_n852,
         mem_stage_inst_dmem_n851, mem_stage_inst_dmem_n850,
         mem_stage_inst_dmem_n849, mem_stage_inst_dmem_n848,
         mem_stage_inst_dmem_n847, mem_stage_inst_dmem_n846,
         mem_stage_inst_dmem_n845, mem_stage_inst_dmem_n844,
         mem_stage_inst_dmem_n843, mem_stage_inst_dmem_n842,
         mem_stage_inst_dmem_n841, mem_stage_inst_dmem_n840,
         mem_stage_inst_dmem_n839, mem_stage_inst_dmem_n838,
         mem_stage_inst_dmem_n837, mem_stage_inst_dmem_n836,
         mem_stage_inst_dmem_n835, mem_stage_inst_dmem_n834,
         mem_stage_inst_dmem_n833, mem_stage_inst_dmem_n832,
         mem_stage_inst_dmem_n831, mem_stage_inst_dmem_n830,
         mem_stage_inst_dmem_n829, mem_stage_inst_dmem_n828,
         mem_stage_inst_dmem_n827, mem_stage_inst_dmem_n826,
         mem_stage_inst_dmem_n825, mem_stage_inst_dmem_n824,
         mem_stage_inst_dmem_n823, mem_stage_inst_dmem_n822,
         mem_stage_inst_dmem_n821, mem_stage_inst_dmem_n820,
         mem_stage_inst_dmem_n819, mem_stage_inst_dmem_n818,
         mem_stage_inst_dmem_n817, mem_stage_inst_dmem_n816,
         mem_stage_inst_dmem_n815, mem_stage_inst_dmem_n814,
         mem_stage_inst_dmem_n813, mem_stage_inst_dmem_n812,
         mem_stage_inst_dmem_n811, mem_stage_inst_dmem_n810,
         mem_stage_inst_dmem_n809, mem_stage_inst_dmem_n808,
         mem_stage_inst_dmem_n807, mem_stage_inst_dmem_n806,
         mem_stage_inst_dmem_n805, mem_stage_inst_dmem_n804,
         mem_stage_inst_dmem_n803, mem_stage_inst_dmem_n802,
         mem_stage_inst_dmem_n801, mem_stage_inst_dmem_n800,
         mem_stage_inst_dmem_n799, mem_stage_inst_dmem_n798,
         mem_stage_inst_dmem_n797, mem_stage_inst_dmem_n796,
         mem_stage_inst_dmem_n795, mem_stage_inst_dmem_n794,
         mem_stage_inst_dmem_n793, mem_stage_inst_dmem_n792,
         mem_stage_inst_dmem_n791, mem_stage_inst_dmem_n790,
         mem_stage_inst_dmem_n789, mem_stage_inst_dmem_n788,
         mem_stage_inst_dmem_n787, mem_stage_inst_dmem_n786,
         mem_stage_inst_dmem_n785, mem_stage_inst_dmem_n784,
         mem_stage_inst_dmem_n783, mem_stage_inst_dmem_n782,
         mem_stage_inst_dmem_n781, mem_stage_inst_dmem_n780,
         mem_stage_inst_dmem_n779, mem_stage_inst_dmem_n778,
         mem_stage_inst_dmem_n777, mem_stage_inst_dmem_n776,
         mem_stage_inst_dmem_n775, mem_stage_inst_dmem_n774,
         mem_stage_inst_dmem_n773, mem_stage_inst_dmem_n772,
         mem_stage_inst_dmem_n771, mem_stage_inst_dmem_n770,
         mem_stage_inst_dmem_n769, mem_stage_inst_dmem_n768,
         mem_stage_inst_dmem_n767, mem_stage_inst_dmem_n766,
         mem_stage_inst_dmem_n765, mem_stage_inst_dmem_n764,
         mem_stage_inst_dmem_n763, mem_stage_inst_dmem_n762,
         mem_stage_inst_dmem_n761, mem_stage_inst_dmem_n760,
         mem_stage_inst_dmem_n759, mem_stage_inst_dmem_n758,
         mem_stage_inst_dmem_n757, mem_stage_inst_dmem_n756,
         mem_stage_inst_dmem_n755, mem_stage_inst_dmem_n754,
         mem_stage_inst_dmem_n753, mem_stage_inst_dmem_n752,
         mem_stage_inst_dmem_n751, mem_stage_inst_dmem_n750,
         mem_stage_inst_dmem_n749, mem_stage_inst_dmem_n748,
         mem_stage_inst_dmem_n747, mem_stage_inst_dmem_n746,
         mem_stage_inst_dmem_n745, mem_stage_inst_dmem_n744,
         mem_stage_inst_dmem_n743, mem_stage_inst_dmem_n742,
         mem_stage_inst_dmem_n741, mem_stage_inst_dmem_n740,
         mem_stage_inst_dmem_n739, mem_stage_inst_dmem_n738,
         mem_stage_inst_dmem_n737, mem_stage_inst_dmem_n736,
         mem_stage_inst_dmem_n735, mem_stage_inst_dmem_n734,
         mem_stage_inst_dmem_n733, mem_stage_inst_dmem_n732,
         mem_stage_inst_dmem_n731, mem_stage_inst_dmem_n730,
         mem_stage_inst_dmem_n729, mem_stage_inst_dmem_n728,
         mem_stage_inst_dmem_n727, mem_stage_inst_dmem_n726,
         mem_stage_inst_dmem_n725, mem_stage_inst_dmem_n724,
         mem_stage_inst_dmem_n723, mem_stage_inst_dmem_n722,
         mem_stage_inst_dmem_n721, mem_stage_inst_dmem_n720,
         mem_stage_inst_dmem_n719, mem_stage_inst_dmem_n718,
         mem_stage_inst_dmem_n717, mem_stage_inst_dmem_n716,
         mem_stage_inst_dmem_n715, mem_stage_inst_dmem_n714,
         mem_stage_inst_dmem_n713, mem_stage_inst_dmem_n712,
         mem_stage_inst_dmem_n711, mem_stage_inst_dmem_n710,
         mem_stage_inst_dmem_n709, mem_stage_inst_dmem_n708,
         mem_stage_inst_dmem_n707, mem_stage_inst_dmem_n706,
         mem_stage_inst_dmem_n705, mem_stage_inst_dmem_n704,
         mem_stage_inst_dmem_n703, mem_stage_inst_dmem_n702,
         mem_stage_inst_dmem_n701, mem_stage_inst_dmem_n700,
         mem_stage_inst_dmem_n699, mem_stage_inst_dmem_n698,
         mem_stage_inst_dmem_n697, mem_stage_inst_dmem_n696,
         mem_stage_inst_dmem_n695, mem_stage_inst_dmem_n694,
         mem_stage_inst_dmem_n693, mem_stage_inst_dmem_n692,
         mem_stage_inst_dmem_n691, mem_stage_inst_dmem_n690,
         mem_stage_inst_dmem_n689, mem_stage_inst_dmem_n688,
         mem_stage_inst_dmem_n687, mem_stage_inst_dmem_n686,
         mem_stage_inst_dmem_n685, mem_stage_inst_dmem_n684,
         mem_stage_inst_dmem_n683, mem_stage_inst_dmem_n682,
         mem_stage_inst_dmem_n681, mem_stage_inst_dmem_n680,
         mem_stage_inst_dmem_n679, mem_stage_inst_dmem_n678,
         mem_stage_inst_dmem_n677, mem_stage_inst_dmem_n676,
         mem_stage_inst_dmem_n675, mem_stage_inst_dmem_n674,
         mem_stage_inst_dmem_n673, mem_stage_inst_dmem_n672,
         mem_stage_inst_dmem_n671, mem_stage_inst_dmem_n670,
         mem_stage_inst_dmem_n669, mem_stage_inst_dmem_n668,
         mem_stage_inst_dmem_n667, mem_stage_inst_dmem_n666,
         mem_stage_inst_dmem_n665, mem_stage_inst_dmem_n664,
         mem_stage_inst_dmem_n663, mem_stage_inst_dmem_n662,
         mem_stage_inst_dmem_n661, mem_stage_inst_dmem_n660,
         mem_stage_inst_dmem_n659, mem_stage_inst_dmem_n658,
         mem_stage_inst_dmem_n657, mem_stage_inst_dmem_n656,
         mem_stage_inst_dmem_n655, mem_stage_inst_dmem_n654,
         mem_stage_inst_dmem_n653, mem_stage_inst_dmem_n652,
         mem_stage_inst_dmem_n651, mem_stage_inst_dmem_n650,
         mem_stage_inst_dmem_n649, mem_stage_inst_dmem_n648,
         mem_stage_inst_dmem_n647, mem_stage_inst_dmem_n646,
         mem_stage_inst_dmem_n645, mem_stage_inst_dmem_n644,
         mem_stage_inst_dmem_n643, mem_stage_inst_dmem_n642,
         mem_stage_inst_dmem_n641, mem_stage_inst_dmem_n640,
         mem_stage_inst_dmem_n639, mem_stage_inst_dmem_n638,
         mem_stage_inst_dmem_n637, mem_stage_inst_dmem_n636,
         mem_stage_inst_dmem_n635, mem_stage_inst_dmem_n634,
         mem_stage_inst_dmem_n633, mem_stage_inst_dmem_n632,
         mem_stage_inst_dmem_n631, mem_stage_inst_dmem_n630,
         mem_stage_inst_dmem_n629, mem_stage_inst_dmem_n628,
         mem_stage_inst_dmem_n627, mem_stage_inst_dmem_n626,
         mem_stage_inst_dmem_n625, mem_stage_inst_dmem_n624,
         mem_stage_inst_dmem_n623, mem_stage_inst_dmem_n622,
         mem_stage_inst_dmem_n621, mem_stage_inst_dmem_n620,
         mem_stage_inst_dmem_n619, mem_stage_inst_dmem_n618,
         mem_stage_inst_dmem_n617, mem_stage_inst_dmem_n616,
         mem_stage_inst_dmem_n615, mem_stage_inst_dmem_n614,
         mem_stage_inst_dmem_n613, mem_stage_inst_dmem_n612,
         mem_stage_inst_dmem_n611, mem_stage_inst_dmem_n610,
         mem_stage_inst_dmem_n609, mem_stage_inst_dmem_n608,
         mem_stage_inst_dmem_n607, mem_stage_inst_dmem_n606,
         mem_stage_inst_dmem_n605, mem_stage_inst_dmem_n604,
         mem_stage_inst_dmem_n603, mem_stage_inst_dmem_n602,
         mem_stage_inst_dmem_n601, mem_stage_inst_dmem_n600,
         mem_stage_inst_dmem_n599, mem_stage_inst_dmem_n598,
         mem_stage_inst_dmem_n597, mem_stage_inst_dmem_n596,
         mem_stage_inst_dmem_n595, mem_stage_inst_dmem_n594,
         mem_stage_inst_dmem_n593, mem_stage_inst_dmem_n592,
         mem_stage_inst_dmem_n591, mem_stage_inst_dmem_n590,
         mem_stage_inst_dmem_n589, mem_stage_inst_dmem_n588,
         mem_stage_inst_dmem_n587, mem_stage_inst_dmem_n586,
         mem_stage_inst_dmem_n585, mem_stage_inst_dmem_n584,
         mem_stage_inst_dmem_n583, mem_stage_inst_dmem_n582,
         mem_stage_inst_dmem_n581, mem_stage_inst_dmem_n580,
         mem_stage_inst_dmem_n579, mem_stage_inst_dmem_n578,
         mem_stage_inst_dmem_n577, mem_stage_inst_dmem_n576,
         mem_stage_inst_dmem_n575, mem_stage_inst_dmem_n574,
         mem_stage_inst_dmem_n573, mem_stage_inst_dmem_n572,
         mem_stage_inst_dmem_n571, mem_stage_inst_dmem_n570,
         mem_stage_inst_dmem_n569, mem_stage_inst_dmem_n568,
         mem_stage_inst_dmem_n567, mem_stage_inst_dmem_n566,
         mem_stage_inst_dmem_n565, mem_stage_inst_dmem_ram_224__0_,
         mem_stage_inst_dmem_ram_224__1_, mem_stage_inst_dmem_ram_224__2_,
         mem_stage_inst_dmem_ram_224__3_, mem_stage_inst_dmem_ram_224__4_,
         mem_stage_inst_dmem_ram_224__5_, mem_stage_inst_dmem_ram_224__6_,
         mem_stage_inst_dmem_ram_224__7_, mem_stage_inst_dmem_ram_224__8_,
         mem_stage_inst_dmem_ram_224__9_, mem_stage_inst_dmem_ram_224__10_,
         mem_stage_inst_dmem_ram_224__11_, mem_stage_inst_dmem_ram_224__12_,
         mem_stage_inst_dmem_ram_224__13_, mem_stage_inst_dmem_ram_224__14_,
         mem_stage_inst_dmem_ram_224__15_, mem_stage_inst_dmem_ram_225__0_,
         mem_stage_inst_dmem_ram_225__1_, mem_stage_inst_dmem_ram_225__2_,
         mem_stage_inst_dmem_ram_225__3_, mem_stage_inst_dmem_ram_225__4_,
         mem_stage_inst_dmem_ram_225__5_, mem_stage_inst_dmem_ram_225__6_,
         mem_stage_inst_dmem_ram_225__7_, mem_stage_inst_dmem_ram_225__8_,
         mem_stage_inst_dmem_ram_225__9_, mem_stage_inst_dmem_ram_225__10_,
         mem_stage_inst_dmem_ram_225__11_, mem_stage_inst_dmem_ram_225__12_,
         mem_stage_inst_dmem_ram_225__13_, mem_stage_inst_dmem_ram_225__14_,
         mem_stage_inst_dmem_ram_225__15_, mem_stage_inst_dmem_ram_226__0_,
         mem_stage_inst_dmem_ram_226__1_, mem_stage_inst_dmem_ram_226__2_,
         mem_stage_inst_dmem_ram_226__3_, mem_stage_inst_dmem_ram_226__4_,
         mem_stage_inst_dmem_ram_226__5_, mem_stage_inst_dmem_ram_226__6_,
         mem_stage_inst_dmem_ram_226__7_, mem_stage_inst_dmem_ram_226__8_,
         mem_stage_inst_dmem_ram_226__9_, mem_stage_inst_dmem_ram_226__10_,
         mem_stage_inst_dmem_ram_226__11_, mem_stage_inst_dmem_ram_226__12_,
         mem_stage_inst_dmem_ram_226__13_, mem_stage_inst_dmem_ram_226__14_,
         mem_stage_inst_dmem_ram_226__15_, mem_stage_inst_dmem_ram_227__0_,
         mem_stage_inst_dmem_ram_227__1_, mem_stage_inst_dmem_ram_227__2_,
         mem_stage_inst_dmem_ram_227__3_, mem_stage_inst_dmem_ram_227__4_,
         mem_stage_inst_dmem_ram_227__5_, mem_stage_inst_dmem_ram_227__6_,
         mem_stage_inst_dmem_ram_227__7_, mem_stage_inst_dmem_ram_227__8_,
         mem_stage_inst_dmem_ram_227__9_, mem_stage_inst_dmem_ram_227__10_,
         mem_stage_inst_dmem_ram_227__11_, mem_stage_inst_dmem_ram_227__12_,
         mem_stage_inst_dmem_ram_227__13_, mem_stage_inst_dmem_ram_227__14_,
         mem_stage_inst_dmem_ram_227__15_, mem_stage_inst_dmem_ram_228__0_,
         mem_stage_inst_dmem_ram_228__1_, mem_stage_inst_dmem_ram_228__2_,
         mem_stage_inst_dmem_ram_228__3_, mem_stage_inst_dmem_ram_228__4_,
         mem_stage_inst_dmem_ram_228__5_, mem_stage_inst_dmem_ram_228__6_,
         mem_stage_inst_dmem_ram_228__7_, mem_stage_inst_dmem_ram_228__8_,
         mem_stage_inst_dmem_ram_228__9_, mem_stage_inst_dmem_ram_228__10_,
         mem_stage_inst_dmem_ram_228__11_, mem_stage_inst_dmem_ram_228__12_,
         mem_stage_inst_dmem_ram_228__13_, mem_stage_inst_dmem_ram_228__14_,
         mem_stage_inst_dmem_ram_228__15_, mem_stage_inst_dmem_ram_229__0_,
         mem_stage_inst_dmem_ram_229__1_, mem_stage_inst_dmem_ram_229__2_,
         mem_stage_inst_dmem_ram_229__3_, mem_stage_inst_dmem_ram_229__4_,
         mem_stage_inst_dmem_ram_229__5_, mem_stage_inst_dmem_ram_229__6_,
         mem_stage_inst_dmem_ram_229__7_, mem_stage_inst_dmem_ram_229__8_,
         mem_stage_inst_dmem_ram_229__9_, mem_stage_inst_dmem_ram_229__10_,
         mem_stage_inst_dmem_ram_229__11_, mem_stage_inst_dmem_ram_229__12_,
         mem_stage_inst_dmem_ram_229__13_, mem_stage_inst_dmem_ram_229__14_,
         mem_stage_inst_dmem_ram_229__15_, mem_stage_inst_dmem_ram_230__0_,
         mem_stage_inst_dmem_ram_230__1_, mem_stage_inst_dmem_ram_230__2_,
         mem_stage_inst_dmem_ram_230__3_, mem_stage_inst_dmem_ram_230__4_,
         mem_stage_inst_dmem_ram_230__5_, mem_stage_inst_dmem_ram_230__6_,
         mem_stage_inst_dmem_ram_230__7_, mem_stage_inst_dmem_ram_230__8_,
         mem_stage_inst_dmem_ram_230__9_, mem_stage_inst_dmem_ram_230__10_,
         mem_stage_inst_dmem_ram_230__11_, mem_stage_inst_dmem_ram_230__12_,
         mem_stage_inst_dmem_ram_230__13_, mem_stage_inst_dmem_ram_230__14_,
         mem_stage_inst_dmem_ram_230__15_, mem_stage_inst_dmem_ram_231__0_,
         mem_stage_inst_dmem_ram_231__1_, mem_stage_inst_dmem_ram_231__2_,
         mem_stage_inst_dmem_ram_231__3_, mem_stage_inst_dmem_ram_231__4_,
         mem_stage_inst_dmem_ram_231__5_, mem_stage_inst_dmem_ram_231__6_,
         mem_stage_inst_dmem_ram_231__7_, mem_stage_inst_dmem_ram_231__8_,
         mem_stage_inst_dmem_ram_231__9_, mem_stage_inst_dmem_ram_231__10_,
         mem_stage_inst_dmem_ram_231__11_, mem_stage_inst_dmem_ram_231__12_,
         mem_stage_inst_dmem_ram_231__13_, mem_stage_inst_dmem_ram_231__14_,
         mem_stage_inst_dmem_ram_231__15_, mem_stage_inst_dmem_ram_232__0_,
         mem_stage_inst_dmem_ram_232__1_, mem_stage_inst_dmem_ram_232__2_,
         mem_stage_inst_dmem_ram_232__3_, mem_stage_inst_dmem_ram_232__4_,
         mem_stage_inst_dmem_ram_232__5_, mem_stage_inst_dmem_ram_232__6_,
         mem_stage_inst_dmem_ram_232__7_, mem_stage_inst_dmem_ram_232__8_,
         mem_stage_inst_dmem_ram_232__9_, mem_stage_inst_dmem_ram_232__10_,
         mem_stage_inst_dmem_ram_232__11_, mem_stage_inst_dmem_ram_232__12_,
         mem_stage_inst_dmem_ram_232__13_, mem_stage_inst_dmem_ram_232__14_,
         mem_stage_inst_dmem_ram_232__15_, mem_stage_inst_dmem_ram_233__0_,
         mem_stage_inst_dmem_ram_233__1_, mem_stage_inst_dmem_ram_233__2_,
         mem_stage_inst_dmem_ram_233__3_, mem_stage_inst_dmem_ram_233__4_,
         mem_stage_inst_dmem_ram_233__5_, mem_stage_inst_dmem_ram_233__6_,
         mem_stage_inst_dmem_ram_233__7_, mem_stage_inst_dmem_ram_233__8_,
         mem_stage_inst_dmem_ram_233__9_, mem_stage_inst_dmem_ram_233__10_,
         mem_stage_inst_dmem_ram_233__11_, mem_stage_inst_dmem_ram_233__12_,
         mem_stage_inst_dmem_ram_233__13_, mem_stage_inst_dmem_ram_233__14_,
         mem_stage_inst_dmem_ram_233__15_, mem_stage_inst_dmem_ram_234__0_,
         mem_stage_inst_dmem_ram_234__1_, mem_stage_inst_dmem_ram_234__2_,
         mem_stage_inst_dmem_ram_234__3_, mem_stage_inst_dmem_ram_234__4_,
         mem_stage_inst_dmem_ram_234__5_, mem_stage_inst_dmem_ram_234__6_,
         mem_stage_inst_dmem_ram_234__7_, mem_stage_inst_dmem_ram_234__8_,
         mem_stage_inst_dmem_ram_234__9_, mem_stage_inst_dmem_ram_234__10_,
         mem_stage_inst_dmem_ram_234__11_, mem_stage_inst_dmem_ram_234__12_,
         mem_stage_inst_dmem_ram_234__13_, mem_stage_inst_dmem_ram_234__14_,
         mem_stage_inst_dmem_ram_234__15_, mem_stage_inst_dmem_ram_235__0_,
         mem_stage_inst_dmem_ram_235__1_, mem_stage_inst_dmem_ram_235__2_,
         mem_stage_inst_dmem_ram_235__3_, mem_stage_inst_dmem_ram_235__4_,
         mem_stage_inst_dmem_ram_235__5_, mem_stage_inst_dmem_ram_235__6_,
         mem_stage_inst_dmem_ram_235__7_, mem_stage_inst_dmem_ram_235__8_,
         mem_stage_inst_dmem_ram_235__9_, mem_stage_inst_dmem_ram_235__10_,
         mem_stage_inst_dmem_ram_235__11_, mem_stage_inst_dmem_ram_235__12_,
         mem_stage_inst_dmem_ram_235__13_, mem_stage_inst_dmem_ram_235__14_,
         mem_stage_inst_dmem_ram_235__15_, mem_stage_inst_dmem_ram_236__0_,
         mem_stage_inst_dmem_ram_236__1_, mem_stage_inst_dmem_ram_236__2_,
         mem_stage_inst_dmem_ram_236__3_, mem_stage_inst_dmem_ram_236__4_,
         mem_stage_inst_dmem_ram_236__5_, mem_stage_inst_dmem_ram_236__6_,
         mem_stage_inst_dmem_ram_236__7_, mem_stage_inst_dmem_ram_236__8_,
         mem_stage_inst_dmem_ram_236__9_, mem_stage_inst_dmem_ram_236__10_,
         mem_stage_inst_dmem_ram_236__11_, mem_stage_inst_dmem_ram_236__12_,
         mem_stage_inst_dmem_ram_236__13_, mem_stage_inst_dmem_ram_236__14_,
         mem_stage_inst_dmem_ram_236__15_, mem_stage_inst_dmem_ram_237__0_,
         mem_stage_inst_dmem_ram_237__1_, mem_stage_inst_dmem_ram_237__2_,
         mem_stage_inst_dmem_ram_237__3_, mem_stage_inst_dmem_ram_237__4_,
         mem_stage_inst_dmem_ram_237__5_, mem_stage_inst_dmem_ram_237__6_,
         mem_stage_inst_dmem_ram_237__7_, mem_stage_inst_dmem_ram_237__8_,
         mem_stage_inst_dmem_ram_237__9_, mem_stage_inst_dmem_ram_237__10_,
         mem_stage_inst_dmem_ram_237__11_, mem_stage_inst_dmem_ram_237__12_,
         mem_stage_inst_dmem_ram_237__13_, mem_stage_inst_dmem_ram_237__14_,
         mem_stage_inst_dmem_ram_237__15_, mem_stage_inst_dmem_ram_238__0_,
         mem_stage_inst_dmem_ram_238__1_, mem_stage_inst_dmem_ram_238__2_,
         mem_stage_inst_dmem_ram_238__3_, mem_stage_inst_dmem_ram_238__4_,
         mem_stage_inst_dmem_ram_238__5_, mem_stage_inst_dmem_ram_238__6_,
         mem_stage_inst_dmem_ram_238__7_, mem_stage_inst_dmem_ram_238__8_,
         mem_stage_inst_dmem_ram_238__9_, mem_stage_inst_dmem_ram_238__10_,
         mem_stage_inst_dmem_ram_238__11_, mem_stage_inst_dmem_ram_238__12_,
         mem_stage_inst_dmem_ram_238__13_, mem_stage_inst_dmem_ram_238__14_,
         mem_stage_inst_dmem_ram_238__15_, mem_stage_inst_dmem_ram_239__0_,
         mem_stage_inst_dmem_ram_239__1_, mem_stage_inst_dmem_ram_239__2_,
         mem_stage_inst_dmem_ram_239__3_, mem_stage_inst_dmem_ram_239__4_,
         mem_stage_inst_dmem_ram_239__5_, mem_stage_inst_dmem_ram_239__6_,
         mem_stage_inst_dmem_ram_239__7_, mem_stage_inst_dmem_ram_239__8_,
         mem_stage_inst_dmem_ram_239__9_, mem_stage_inst_dmem_ram_239__10_,
         mem_stage_inst_dmem_ram_239__11_, mem_stage_inst_dmem_ram_239__12_,
         mem_stage_inst_dmem_ram_239__13_, mem_stage_inst_dmem_ram_239__14_,
         mem_stage_inst_dmem_ram_239__15_, mem_stage_inst_dmem_ram_240__0_,
         mem_stage_inst_dmem_ram_240__1_, mem_stage_inst_dmem_ram_240__2_,
         mem_stage_inst_dmem_ram_240__3_, mem_stage_inst_dmem_ram_240__4_,
         mem_stage_inst_dmem_ram_240__5_, mem_stage_inst_dmem_ram_240__6_,
         mem_stage_inst_dmem_ram_240__7_, mem_stage_inst_dmem_ram_240__8_,
         mem_stage_inst_dmem_ram_240__9_, mem_stage_inst_dmem_ram_240__10_,
         mem_stage_inst_dmem_ram_240__11_, mem_stage_inst_dmem_ram_240__12_,
         mem_stage_inst_dmem_ram_240__13_, mem_stage_inst_dmem_ram_240__14_,
         mem_stage_inst_dmem_ram_240__15_, mem_stage_inst_dmem_ram_241__0_,
         mem_stage_inst_dmem_ram_241__1_, mem_stage_inst_dmem_ram_241__2_,
         mem_stage_inst_dmem_ram_241__3_, mem_stage_inst_dmem_ram_241__4_,
         mem_stage_inst_dmem_ram_241__5_, mem_stage_inst_dmem_ram_241__6_,
         mem_stage_inst_dmem_ram_241__7_, mem_stage_inst_dmem_ram_241__8_,
         mem_stage_inst_dmem_ram_241__9_, mem_stage_inst_dmem_ram_241__10_,
         mem_stage_inst_dmem_ram_241__11_, mem_stage_inst_dmem_ram_241__12_,
         mem_stage_inst_dmem_ram_241__13_, mem_stage_inst_dmem_ram_241__14_,
         mem_stage_inst_dmem_ram_241__15_, mem_stage_inst_dmem_ram_242__0_,
         mem_stage_inst_dmem_ram_242__1_, mem_stage_inst_dmem_ram_242__2_,
         mem_stage_inst_dmem_ram_242__3_, mem_stage_inst_dmem_ram_242__4_,
         mem_stage_inst_dmem_ram_242__5_, mem_stage_inst_dmem_ram_242__6_,
         mem_stage_inst_dmem_ram_242__7_, mem_stage_inst_dmem_ram_242__8_,
         mem_stage_inst_dmem_ram_242__9_, mem_stage_inst_dmem_ram_242__10_,
         mem_stage_inst_dmem_ram_242__11_, mem_stage_inst_dmem_ram_242__12_,
         mem_stage_inst_dmem_ram_242__13_, mem_stage_inst_dmem_ram_242__14_,
         mem_stage_inst_dmem_ram_242__15_, mem_stage_inst_dmem_ram_243__0_,
         mem_stage_inst_dmem_ram_243__1_, mem_stage_inst_dmem_ram_243__2_,
         mem_stage_inst_dmem_ram_243__3_, mem_stage_inst_dmem_ram_243__4_,
         mem_stage_inst_dmem_ram_243__5_, mem_stage_inst_dmem_ram_243__6_,
         mem_stage_inst_dmem_ram_243__7_, mem_stage_inst_dmem_ram_243__8_,
         mem_stage_inst_dmem_ram_243__9_, mem_stage_inst_dmem_ram_243__10_,
         mem_stage_inst_dmem_ram_243__11_, mem_stage_inst_dmem_ram_243__12_,
         mem_stage_inst_dmem_ram_243__13_, mem_stage_inst_dmem_ram_243__14_,
         mem_stage_inst_dmem_ram_243__15_, mem_stage_inst_dmem_ram_244__0_,
         mem_stage_inst_dmem_ram_244__1_, mem_stage_inst_dmem_ram_244__2_,
         mem_stage_inst_dmem_ram_244__3_, mem_stage_inst_dmem_ram_244__4_,
         mem_stage_inst_dmem_ram_244__5_, mem_stage_inst_dmem_ram_244__6_,
         mem_stage_inst_dmem_ram_244__7_, mem_stage_inst_dmem_ram_244__8_,
         mem_stage_inst_dmem_ram_244__9_, mem_stage_inst_dmem_ram_244__10_,
         mem_stage_inst_dmem_ram_244__11_, mem_stage_inst_dmem_ram_244__12_,
         mem_stage_inst_dmem_ram_244__13_, mem_stage_inst_dmem_ram_244__14_,
         mem_stage_inst_dmem_ram_244__15_, mem_stage_inst_dmem_ram_245__0_,
         mem_stage_inst_dmem_ram_245__1_, mem_stage_inst_dmem_ram_245__2_,
         mem_stage_inst_dmem_ram_245__3_, mem_stage_inst_dmem_ram_245__4_,
         mem_stage_inst_dmem_ram_245__5_, mem_stage_inst_dmem_ram_245__6_,
         mem_stage_inst_dmem_ram_245__7_, mem_stage_inst_dmem_ram_245__8_,
         mem_stage_inst_dmem_ram_245__9_, mem_stage_inst_dmem_ram_245__10_,
         mem_stage_inst_dmem_ram_245__11_, mem_stage_inst_dmem_ram_245__12_,
         mem_stage_inst_dmem_ram_245__13_, mem_stage_inst_dmem_ram_245__14_,
         mem_stage_inst_dmem_ram_245__15_, mem_stage_inst_dmem_ram_246__0_,
         mem_stage_inst_dmem_ram_246__1_, mem_stage_inst_dmem_ram_246__2_,
         mem_stage_inst_dmem_ram_246__3_, mem_stage_inst_dmem_ram_246__4_,
         mem_stage_inst_dmem_ram_246__5_, mem_stage_inst_dmem_ram_246__6_,
         mem_stage_inst_dmem_ram_246__7_, mem_stage_inst_dmem_ram_246__8_,
         mem_stage_inst_dmem_ram_246__9_, mem_stage_inst_dmem_ram_246__10_,
         mem_stage_inst_dmem_ram_246__11_, mem_stage_inst_dmem_ram_246__12_,
         mem_stage_inst_dmem_ram_246__13_, mem_stage_inst_dmem_ram_246__14_,
         mem_stage_inst_dmem_ram_246__15_, mem_stage_inst_dmem_ram_247__0_,
         mem_stage_inst_dmem_ram_247__1_, mem_stage_inst_dmem_ram_247__2_,
         mem_stage_inst_dmem_ram_247__3_, mem_stage_inst_dmem_ram_247__4_,
         mem_stage_inst_dmem_ram_247__5_, mem_stage_inst_dmem_ram_247__6_,
         mem_stage_inst_dmem_ram_247__7_, mem_stage_inst_dmem_ram_247__8_,
         mem_stage_inst_dmem_ram_247__9_, mem_stage_inst_dmem_ram_247__10_,
         mem_stage_inst_dmem_ram_247__11_, mem_stage_inst_dmem_ram_247__12_,
         mem_stage_inst_dmem_ram_247__13_, mem_stage_inst_dmem_ram_247__14_,
         mem_stage_inst_dmem_ram_247__15_, mem_stage_inst_dmem_ram_248__0_,
         mem_stage_inst_dmem_ram_248__1_, mem_stage_inst_dmem_ram_248__2_,
         mem_stage_inst_dmem_ram_248__3_, mem_stage_inst_dmem_ram_248__4_,
         mem_stage_inst_dmem_ram_248__5_, mem_stage_inst_dmem_ram_248__6_,
         mem_stage_inst_dmem_ram_248__7_, mem_stage_inst_dmem_ram_248__8_,
         mem_stage_inst_dmem_ram_248__9_, mem_stage_inst_dmem_ram_248__10_,
         mem_stage_inst_dmem_ram_248__11_, mem_stage_inst_dmem_ram_248__12_,
         mem_stage_inst_dmem_ram_248__13_, mem_stage_inst_dmem_ram_248__14_,
         mem_stage_inst_dmem_ram_248__15_, mem_stage_inst_dmem_ram_249__0_,
         mem_stage_inst_dmem_ram_249__1_, mem_stage_inst_dmem_ram_249__2_,
         mem_stage_inst_dmem_ram_249__3_, mem_stage_inst_dmem_ram_249__4_,
         mem_stage_inst_dmem_ram_249__5_, mem_stage_inst_dmem_ram_249__6_,
         mem_stage_inst_dmem_ram_249__7_, mem_stage_inst_dmem_ram_249__8_,
         mem_stage_inst_dmem_ram_249__9_, mem_stage_inst_dmem_ram_249__10_,
         mem_stage_inst_dmem_ram_249__11_, mem_stage_inst_dmem_ram_249__12_,
         mem_stage_inst_dmem_ram_249__13_, mem_stage_inst_dmem_ram_249__14_,
         mem_stage_inst_dmem_ram_249__15_, mem_stage_inst_dmem_ram_250__0_,
         mem_stage_inst_dmem_ram_250__1_, mem_stage_inst_dmem_ram_250__2_,
         mem_stage_inst_dmem_ram_250__3_, mem_stage_inst_dmem_ram_250__4_,
         mem_stage_inst_dmem_ram_250__5_, mem_stage_inst_dmem_ram_250__6_,
         mem_stage_inst_dmem_ram_250__7_, mem_stage_inst_dmem_ram_250__8_,
         mem_stage_inst_dmem_ram_250__9_, mem_stage_inst_dmem_ram_250__10_,
         mem_stage_inst_dmem_ram_250__11_, mem_stage_inst_dmem_ram_250__12_,
         mem_stage_inst_dmem_ram_250__13_, mem_stage_inst_dmem_ram_250__14_,
         mem_stage_inst_dmem_ram_250__15_, mem_stage_inst_dmem_ram_251__0_,
         mem_stage_inst_dmem_ram_251__1_, mem_stage_inst_dmem_ram_251__2_,
         mem_stage_inst_dmem_ram_251__3_, mem_stage_inst_dmem_ram_251__4_,
         mem_stage_inst_dmem_ram_251__5_, mem_stage_inst_dmem_ram_251__6_,
         mem_stage_inst_dmem_ram_251__7_, mem_stage_inst_dmem_ram_251__8_,
         mem_stage_inst_dmem_ram_251__9_, mem_stage_inst_dmem_ram_251__10_,
         mem_stage_inst_dmem_ram_251__11_, mem_stage_inst_dmem_ram_251__12_,
         mem_stage_inst_dmem_ram_251__13_, mem_stage_inst_dmem_ram_251__14_,
         mem_stage_inst_dmem_ram_251__15_, mem_stage_inst_dmem_ram_252__0_,
         mem_stage_inst_dmem_ram_252__1_, mem_stage_inst_dmem_ram_252__2_,
         mem_stage_inst_dmem_ram_252__3_, mem_stage_inst_dmem_ram_252__4_,
         mem_stage_inst_dmem_ram_252__5_, mem_stage_inst_dmem_ram_252__6_,
         mem_stage_inst_dmem_ram_252__7_, mem_stage_inst_dmem_ram_252__8_,
         mem_stage_inst_dmem_ram_252__9_, mem_stage_inst_dmem_ram_252__10_,
         mem_stage_inst_dmem_ram_252__11_, mem_stage_inst_dmem_ram_252__12_,
         mem_stage_inst_dmem_ram_252__13_, mem_stage_inst_dmem_ram_252__14_,
         mem_stage_inst_dmem_ram_252__15_, mem_stage_inst_dmem_ram_253__0_,
         mem_stage_inst_dmem_ram_253__1_, mem_stage_inst_dmem_ram_253__2_,
         mem_stage_inst_dmem_ram_253__3_, mem_stage_inst_dmem_ram_253__4_,
         mem_stage_inst_dmem_ram_253__5_, mem_stage_inst_dmem_ram_253__6_,
         mem_stage_inst_dmem_ram_253__7_, mem_stage_inst_dmem_ram_253__8_,
         mem_stage_inst_dmem_ram_253__9_, mem_stage_inst_dmem_ram_253__10_,
         mem_stage_inst_dmem_ram_253__11_, mem_stage_inst_dmem_ram_253__12_,
         mem_stage_inst_dmem_ram_253__13_, mem_stage_inst_dmem_ram_253__14_,
         mem_stage_inst_dmem_ram_253__15_, mem_stage_inst_dmem_ram_254__0_,
         mem_stage_inst_dmem_ram_254__1_, mem_stage_inst_dmem_ram_254__2_,
         mem_stage_inst_dmem_ram_254__3_, mem_stage_inst_dmem_ram_254__4_,
         mem_stage_inst_dmem_ram_254__5_, mem_stage_inst_dmem_ram_254__6_,
         mem_stage_inst_dmem_ram_254__7_, mem_stage_inst_dmem_ram_254__8_,
         mem_stage_inst_dmem_ram_254__9_, mem_stage_inst_dmem_ram_254__10_,
         mem_stage_inst_dmem_ram_254__11_, mem_stage_inst_dmem_ram_254__12_,
         mem_stage_inst_dmem_ram_254__13_, mem_stage_inst_dmem_ram_254__14_,
         mem_stage_inst_dmem_ram_254__15_, mem_stage_inst_dmem_ram_255__0_,
         mem_stage_inst_dmem_ram_255__1_, mem_stage_inst_dmem_ram_255__2_,
         mem_stage_inst_dmem_ram_255__3_, mem_stage_inst_dmem_ram_255__4_,
         mem_stage_inst_dmem_ram_255__5_, mem_stage_inst_dmem_ram_255__6_,
         mem_stage_inst_dmem_ram_255__7_, mem_stage_inst_dmem_ram_255__8_,
         mem_stage_inst_dmem_ram_255__9_, mem_stage_inst_dmem_ram_255__10_,
         mem_stage_inst_dmem_ram_255__11_, mem_stage_inst_dmem_ram_255__12_,
         mem_stage_inst_dmem_ram_255__13_, mem_stage_inst_dmem_ram_255__14_,
         mem_stage_inst_dmem_ram_255__15_, mem_stage_inst_dmem_ram_192__0_,
         mem_stage_inst_dmem_ram_192__1_, mem_stage_inst_dmem_ram_192__2_,
         mem_stage_inst_dmem_ram_192__3_, mem_stage_inst_dmem_ram_192__4_,
         mem_stage_inst_dmem_ram_192__5_, mem_stage_inst_dmem_ram_192__6_,
         mem_stage_inst_dmem_ram_192__7_, mem_stage_inst_dmem_ram_192__8_,
         mem_stage_inst_dmem_ram_192__9_, mem_stage_inst_dmem_ram_192__10_,
         mem_stage_inst_dmem_ram_192__11_, mem_stage_inst_dmem_ram_192__12_,
         mem_stage_inst_dmem_ram_192__13_, mem_stage_inst_dmem_ram_192__14_,
         mem_stage_inst_dmem_ram_192__15_, mem_stage_inst_dmem_ram_193__0_,
         mem_stage_inst_dmem_ram_193__1_, mem_stage_inst_dmem_ram_193__2_,
         mem_stage_inst_dmem_ram_193__3_, mem_stage_inst_dmem_ram_193__4_,
         mem_stage_inst_dmem_ram_193__5_, mem_stage_inst_dmem_ram_193__6_,
         mem_stage_inst_dmem_ram_193__7_, mem_stage_inst_dmem_ram_193__8_,
         mem_stage_inst_dmem_ram_193__9_, mem_stage_inst_dmem_ram_193__10_,
         mem_stage_inst_dmem_ram_193__11_, mem_stage_inst_dmem_ram_193__12_,
         mem_stage_inst_dmem_ram_193__13_, mem_stage_inst_dmem_ram_193__14_,
         mem_stage_inst_dmem_ram_193__15_, mem_stage_inst_dmem_ram_194__0_,
         mem_stage_inst_dmem_ram_194__1_, mem_stage_inst_dmem_ram_194__2_,
         mem_stage_inst_dmem_ram_194__3_, mem_stage_inst_dmem_ram_194__4_,
         mem_stage_inst_dmem_ram_194__5_, mem_stage_inst_dmem_ram_194__6_,
         mem_stage_inst_dmem_ram_194__7_, mem_stage_inst_dmem_ram_194__8_,
         mem_stage_inst_dmem_ram_194__9_, mem_stage_inst_dmem_ram_194__10_,
         mem_stage_inst_dmem_ram_194__11_, mem_stage_inst_dmem_ram_194__12_,
         mem_stage_inst_dmem_ram_194__13_, mem_stage_inst_dmem_ram_194__14_,
         mem_stage_inst_dmem_ram_194__15_, mem_stage_inst_dmem_ram_195__0_,
         mem_stage_inst_dmem_ram_195__1_, mem_stage_inst_dmem_ram_195__2_,
         mem_stage_inst_dmem_ram_195__3_, mem_stage_inst_dmem_ram_195__4_,
         mem_stage_inst_dmem_ram_195__5_, mem_stage_inst_dmem_ram_195__6_,
         mem_stage_inst_dmem_ram_195__7_, mem_stage_inst_dmem_ram_195__8_,
         mem_stage_inst_dmem_ram_195__9_, mem_stage_inst_dmem_ram_195__10_,
         mem_stage_inst_dmem_ram_195__11_, mem_stage_inst_dmem_ram_195__12_,
         mem_stage_inst_dmem_ram_195__13_, mem_stage_inst_dmem_ram_195__14_,
         mem_stage_inst_dmem_ram_195__15_, mem_stage_inst_dmem_ram_196__0_,
         mem_stage_inst_dmem_ram_196__1_, mem_stage_inst_dmem_ram_196__2_,
         mem_stage_inst_dmem_ram_196__3_, mem_stage_inst_dmem_ram_196__4_,
         mem_stage_inst_dmem_ram_196__5_, mem_stage_inst_dmem_ram_196__6_,
         mem_stage_inst_dmem_ram_196__7_, mem_stage_inst_dmem_ram_196__8_,
         mem_stage_inst_dmem_ram_196__9_, mem_stage_inst_dmem_ram_196__10_,
         mem_stage_inst_dmem_ram_196__11_, mem_stage_inst_dmem_ram_196__12_,
         mem_stage_inst_dmem_ram_196__13_, mem_stage_inst_dmem_ram_196__14_,
         mem_stage_inst_dmem_ram_196__15_, mem_stage_inst_dmem_ram_197__0_,
         mem_stage_inst_dmem_ram_197__1_, mem_stage_inst_dmem_ram_197__2_,
         mem_stage_inst_dmem_ram_197__3_, mem_stage_inst_dmem_ram_197__4_,
         mem_stage_inst_dmem_ram_197__5_, mem_stage_inst_dmem_ram_197__6_,
         mem_stage_inst_dmem_ram_197__7_, mem_stage_inst_dmem_ram_197__8_,
         mem_stage_inst_dmem_ram_197__9_, mem_stage_inst_dmem_ram_197__10_,
         mem_stage_inst_dmem_ram_197__11_, mem_stage_inst_dmem_ram_197__12_,
         mem_stage_inst_dmem_ram_197__13_, mem_stage_inst_dmem_ram_197__14_,
         mem_stage_inst_dmem_ram_197__15_, mem_stage_inst_dmem_ram_198__0_,
         mem_stage_inst_dmem_ram_198__1_, mem_stage_inst_dmem_ram_198__2_,
         mem_stage_inst_dmem_ram_198__3_, mem_stage_inst_dmem_ram_198__4_,
         mem_stage_inst_dmem_ram_198__5_, mem_stage_inst_dmem_ram_198__6_,
         mem_stage_inst_dmem_ram_198__7_, mem_stage_inst_dmem_ram_198__8_,
         mem_stage_inst_dmem_ram_198__9_, mem_stage_inst_dmem_ram_198__10_,
         mem_stage_inst_dmem_ram_198__11_, mem_stage_inst_dmem_ram_198__12_,
         mem_stage_inst_dmem_ram_198__13_, mem_stage_inst_dmem_ram_198__14_,
         mem_stage_inst_dmem_ram_198__15_, mem_stage_inst_dmem_ram_199__0_,
         mem_stage_inst_dmem_ram_199__1_, mem_stage_inst_dmem_ram_199__2_,
         mem_stage_inst_dmem_ram_199__3_, mem_stage_inst_dmem_ram_199__4_,
         mem_stage_inst_dmem_ram_199__5_, mem_stage_inst_dmem_ram_199__6_,
         mem_stage_inst_dmem_ram_199__7_, mem_stage_inst_dmem_ram_199__8_,
         mem_stage_inst_dmem_ram_199__9_, mem_stage_inst_dmem_ram_199__10_,
         mem_stage_inst_dmem_ram_199__11_, mem_stage_inst_dmem_ram_199__12_,
         mem_stage_inst_dmem_ram_199__13_, mem_stage_inst_dmem_ram_199__14_,
         mem_stage_inst_dmem_ram_199__15_, mem_stage_inst_dmem_ram_200__0_,
         mem_stage_inst_dmem_ram_200__1_, mem_stage_inst_dmem_ram_200__2_,
         mem_stage_inst_dmem_ram_200__3_, mem_stage_inst_dmem_ram_200__4_,
         mem_stage_inst_dmem_ram_200__5_, mem_stage_inst_dmem_ram_200__6_,
         mem_stage_inst_dmem_ram_200__7_, mem_stage_inst_dmem_ram_200__8_,
         mem_stage_inst_dmem_ram_200__9_, mem_stage_inst_dmem_ram_200__10_,
         mem_stage_inst_dmem_ram_200__11_, mem_stage_inst_dmem_ram_200__12_,
         mem_stage_inst_dmem_ram_200__13_, mem_stage_inst_dmem_ram_200__14_,
         mem_stage_inst_dmem_ram_200__15_, mem_stage_inst_dmem_ram_201__0_,
         mem_stage_inst_dmem_ram_201__1_, mem_stage_inst_dmem_ram_201__2_,
         mem_stage_inst_dmem_ram_201__3_, mem_stage_inst_dmem_ram_201__4_,
         mem_stage_inst_dmem_ram_201__5_, mem_stage_inst_dmem_ram_201__6_,
         mem_stage_inst_dmem_ram_201__7_, mem_stage_inst_dmem_ram_201__8_,
         mem_stage_inst_dmem_ram_201__9_, mem_stage_inst_dmem_ram_201__10_,
         mem_stage_inst_dmem_ram_201__11_, mem_stage_inst_dmem_ram_201__12_,
         mem_stage_inst_dmem_ram_201__13_, mem_stage_inst_dmem_ram_201__14_,
         mem_stage_inst_dmem_ram_201__15_, mem_stage_inst_dmem_ram_202__0_,
         mem_stage_inst_dmem_ram_202__1_, mem_stage_inst_dmem_ram_202__2_,
         mem_stage_inst_dmem_ram_202__3_, mem_stage_inst_dmem_ram_202__4_,
         mem_stage_inst_dmem_ram_202__5_, mem_stage_inst_dmem_ram_202__6_,
         mem_stage_inst_dmem_ram_202__7_, mem_stage_inst_dmem_ram_202__8_,
         mem_stage_inst_dmem_ram_202__9_, mem_stage_inst_dmem_ram_202__10_,
         mem_stage_inst_dmem_ram_202__11_, mem_stage_inst_dmem_ram_202__12_,
         mem_stage_inst_dmem_ram_202__13_, mem_stage_inst_dmem_ram_202__14_,
         mem_stage_inst_dmem_ram_202__15_, mem_stage_inst_dmem_ram_203__0_,
         mem_stage_inst_dmem_ram_203__1_, mem_stage_inst_dmem_ram_203__2_,
         mem_stage_inst_dmem_ram_203__3_, mem_stage_inst_dmem_ram_203__4_,
         mem_stage_inst_dmem_ram_203__5_, mem_stage_inst_dmem_ram_203__6_,
         mem_stage_inst_dmem_ram_203__7_, mem_stage_inst_dmem_ram_203__8_,
         mem_stage_inst_dmem_ram_203__9_, mem_stage_inst_dmem_ram_203__10_,
         mem_stage_inst_dmem_ram_203__11_, mem_stage_inst_dmem_ram_203__12_,
         mem_stage_inst_dmem_ram_203__13_, mem_stage_inst_dmem_ram_203__14_,
         mem_stage_inst_dmem_ram_203__15_, mem_stage_inst_dmem_ram_204__0_,
         mem_stage_inst_dmem_ram_204__1_, mem_stage_inst_dmem_ram_204__2_,
         mem_stage_inst_dmem_ram_204__3_, mem_stage_inst_dmem_ram_204__4_,
         mem_stage_inst_dmem_ram_204__5_, mem_stage_inst_dmem_ram_204__6_,
         mem_stage_inst_dmem_ram_204__7_, mem_stage_inst_dmem_ram_204__8_,
         mem_stage_inst_dmem_ram_204__9_, mem_stage_inst_dmem_ram_204__10_,
         mem_stage_inst_dmem_ram_204__11_, mem_stage_inst_dmem_ram_204__12_,
         mem_stage_inst_dmem_ram_204__13_, mem_stage_inst_dmem_ram_204__14_,
         mem_stage_inst_dmem_ram_204__15_, mem_stage_inst_dmem_ram_205__0_,
         mem_stage_inst_dmem_ram_205__1_, mem_stage_inst_dmem_ram_205__2_,
         mem_stage_inst_dmem_ram_205__3_, mem_stage_inst_dmem_ram_205__4_,
         mem_stage_inst_dmem_ram_205__5_, mem_stage_inst_dmem_ram_205__6_,
         mem_stage_inst_dmem_ram_205__7_, mem_stage_inst_dmem_ram_205__8_,
         mem_stage_inst_dmem_ram_205__9_, mem_stage_inst_dmem_ram_205__10_,
         mem_stage_inst_dmem_ram_205__11_, mem_stage_inst_dmem_ram_205__12_,
         mem_stage_inst_dmem_ram_205__13_, mem_stage_inst_dmem_ram_205__14_,
         mem_stage_inst_dmem_ram_205__15_, mem_stage_inst_dmem_ram_206__0_,
         mem_stage_inst_dmem_ram_206__1_, mem_stage_inst_dmem_ram_206__2_,
         mem_stage_inst_dmem_ram_206__3_, mem_stage_inst_dmem_ram_206__4_,
         mem_stage_inst_dmem_ram_206__5_, mem_stage_inst_dmem_ram_206__6_,
         mem_stage_inst_dmem_ram_206__7_, mem_stage_inst_dmem_ram_206__8_,
         mem_stage_inst_dmem_ram_206__9_, mem_stage_inst_dmem_ram_206__10_,
         mem_stage_inst_dmem_ram_206__11_, mem_stage_inst_dmem_ram_206__12_,
         mem_stage_inst_dmem_ram_206__13_, mem_stage_inst_dmem_ram_206__14_,
         mem_stage_inst_dmem_ram_206__15_, mem_stage_inst_dmem_ram_207__0_,
         mem_stage_inst_dmem_ram_207__1_, mem_stage_inst_dmem_ram_207__2_,
         mem_stage_inst_dmem_ram_207__3_, mem_stage_inst_dmem_ram_207__4_,
         mem_stage_inst_dmem_ram_207__5_, mem_stage_inst_dmem_ram_207__6_,
         mem_stage_inst_dmem_ram_207__7_, mem_stage_inst_dmem_ram_207__8_,
         mem_stage_inst_dmem_ram_207__9_, mem_stage_inst_dmem_ram_207__10_,
         mem_stage_inst_dmem_ram_207__11_, mem_stage_inst_dmem_ram_207__12_,
         mem_stage_inst_dmem_ram_207__13_, mem_stage_inst_dmem_ram_207__14_,
         mem_stage_inst_dmem_ram_207__15_, mem_stage_inst_dmem_ram_208__0_,
         mem_stage_inst_dmem_ram_208__1_, mem_stage_inst_dmem_ram_208__2_,
         mem_stage_inst_dmem_ram_208__3_, mem_stage_inst_dmem_ram_208__4_,
         mem_stage_inst_dmem_ram_208__5_, mem_stage_inst_dmem_ram_208__6_,
         mem_stage_inst_dmem_ram_208__7_, mem_stage_inst_dmem_ram_208__8_,
         mem_stage_inst_dmem_ram_208__9_, mem_stage_inst_dmem_ram_208__10_,
         mem_stage_inst_dmem_ram_208__11_, mem_stage_inst_dmem_ram_208__12_,
         mem_stage_inst_dmem_ram_208__13_, mem_stage_inst_dmem_ram_208__14_,
         mem_stage_inst_dmem_ram_208__15_, mem_stage_inst_dmem_ram_209__0_,
         mem_stage_inst_dmem_ram_209__1_, mem_stage_inst_dmem_ram_209__2_,
         mem_stage_inst_dmem_ram_209__3_, mem_stage_inst_dmem_ram_209__4_,
         mem_stage_inst_dmem_ram_209__5_, mem_stage_inst_dmem_ram_209__6_,
         mem_stage_inst_dmem_ram_209__7_, mem_stage_inst_dmem_ram_209__8_,
         mem_stage_inst_dmem_ram_209__9_, mem_stage_inst_dmem_ram_209__10_,
         mem_stage_inst_dmem_ram_209__11_, mem_stage_inst_dmem_ram_209__12_,
         mem_stage_inst_dmem_ram_209__13_, mem_stage_inst_dmem_ram_209__14_,
         mem_stage_inst_dmem_ram_209__15_, mem_stage_inst_dmem_ram_210__0_,
         mem_stage_inst_dmem_ram_210__1_, mem_stage_inst_dmem_ram_210__2_,
         mem_stage_inst_dmem_ram_210__3_, mem_stage_inst_dmem_ram_210__4_,
         mem_stage_inst_dmem_ram_210__5_, mem_stage_inst_dmem_ram_210__6_,
         mem_stage_inst_dmem_ram_210__7_, mem_stage_inst_dmem_ram_210__8_,
         mem_stage_inst_dmem_ram_210__9_, mem_stage_inst_dmem_ram_210__10_,
         mem_stage_inst_dmem_ram_210__11_, mem_stage_inst_dmem_ram_210__12_,
         mem_stage_inst_dmem_ram_210__13_, mem_stage_inst_dmem_ram_210__14_,
         mem_stage_inst_dmem_ram_210__15_, mem_stage_inst_dmem_ram_211__0_,
         mem_stage_inst_dmem_ram_211__1_, mem_stage_inst_dmem_ram_211__2_,
         mem_stage_inst_dmem_ram_211__3_, mem_stage_inst_dmem_ram_211__4_,
         mem_stage_inst_dmem_ram_211__5_, mem_stage_inst_dmem_ram_211__6_,
         mem_stage_inst_dmem_ram_211__7_, mem_stage_inst_dmem_ram_211__8_,
         mem_stage_inst_dmem_ram_211__9_, mem_stage_inst_dmem_ram_211__10_,
         mem_stage_inst_dmem_ram_211__11_, mem_stage_inst_dmem_ram_211__12_,
         mem_stage_inst_dmem_ram_211__13_, mem_stage_inst_dmem_ram_211__14_,
         mem_stage_inst_dmem_ram_211__15_, mem_stage_inst_dmem_ram_212__0_,
         mem_stage_inst_dmem_ram_212__1_, mem_stage_inst_dmem_ram_212__2_,
         mem_stage_inst_dmem_ram_212__3_, mem_stage_inst_dmem_ram_212__4_,
         mem_stage_inst_dmem_ram_212__5_, mem_stage_inst_dmem_ram_212__6_,
         mem_stage_inst_dmem_ram_212__7_, mem_stage_inst_dmem_ram_212__8_,
         mem_stage_inst_dmem_ram_212__9_, mem_stage_inst_dmem_ram_212__10_,
         mem_stage_inst_dmem_ram_212__11_, mem_stage_inst_dmem_ram_212__12_,
         mem_stage_inst_dmem_ram_212__13_, mem_stage_inst_dmem_ram_212__14_,
         mem_stage_inst_dmem_ram_212__15_, mem_stage_inst_dmem_ram_213__0_,
         mem_stage_inst_dmem_ram_213__1_, mem_stage_inst_dmem_ram_213__2_,
         mem_stage_inst_dmem_ram_213__3_, mem_stage_inst_dmem_ram_213__4_,
         mem_stage_inst_dmem_ram_213__5_, mem_stage_inst_dmem_ram_213__6_,
         mem_stage_inst_dmem_ram_213__7_, mem_stage_inst_dmem_ram_213__8_,
         mem_stage_inst_dmem_ram_213__9_, mem_stage_inst_dmem_ram_213__10_,
         mem_stage_inst_dmem_ram_213__11_, mem_stage_inst_dmem_ram_213__12_,
         mem_stage_inst_dmem_ram_213__13_, mem_stage_inst_dmem_ram_213__14_,
         mem_stage_inst_dmem_ram_213__15_, mem_stage_inst_dmem_ram_214__0_,
         mem_stage_inst_dmem_ram_214__1_, mem_stage_inst_dmem_ram_214__2_,
         mem_stage_inst_dmem_ram_214__3_, mem_stage_inst_dmem_ram_214__4_,
         mem_stage_inst_dmem_ram_214__5_, mem_stage_inst_dmem_ram_214__6_,
         mem_stage_inst_dmem_ram_214__7_, mem_stage_inst_dmem_ram_214__8_,
         mem_stage_inst_dmem_ram_214__9_, mem_stage_inst_dmem_ram_214__10_,
         mem_stage_inst_dmem_ram_214__11_, mem_stage_inst_dmem_ram_214__12_,
         mem_stage_inst_dmem_ram_214__13_, mem_stage_inst_dmem_ram_214__14_,
         mem_stage_inst_dmem_ram_214__15_, mem_stage_inst_dmem_ram_215__0_,
         mem_stage_inst_dmem_ram_215__1_, mem_stage_inst_dmem_ram_215__2_,
         mem_stage_inst_dmem_ram_215__3_, mem_stage_inst_dmem_ram_215__4_,
         mem_stage_inst_dmem_ram_215__5_, mem_stage_inst_dmem_ram_215__6_,
         mem_stage_inst_dmem_ram_215__7_, mem_stage_inst_dmem_ram_215__8_,
         mem_stage_inst_dmem_ram_215__9_, mem_stage_inst_dmem_ram_215__10_,
         mem_stage_inst_dmem_ram_215__11_, mem_stage_inst_dmem_ram_215__12_,
         mem_stage_inst_dmem_ram_215__13_, mem_stage_inst_dmem_ram_215__14_,
         mem_stage_inst_dmem_ram_215__15_, mem_stage_inst_dmem_ram_216__0_,
         mem_stage_inst_dmem_ram_216__1_, mem_stage_inst_dmem_ram_216__2_,
         mem_stage_inst_dmem_ram_216__3_, mem_stage_inst_dmem_ram_216__4_,
         mem_stage_inst_dmem_ram_216__5_, mem_stage_inst_dmem_ram_216__6_,
         mem_stage_inst_dmem_ram_216__7_, mem_stage_inst_dmem_ram_216__8_,
         mem_stage_inst_dmem_ram_216__9_, mem_stage_inst_dmem_ram_216__10_,
         mem_stage_inst_dmem_ram_216__11_, mem_stage_inst_dmem_ram_216__12_,
         mem_stage_inst_dmem_ram_216__13_, mem_stage_inst_dmem_ram_216__14_,
         mem_stage_inst_dmem_ram_216__15_, mem_stage_inst_dmem_ram_217__0_,
         mem_stage_inst_dmem_ram_217__1_, mem_stage_inst_dmem_ram_217__2_,
         mem_stage_inst_dmem_ram_217__3_, mem_stage_inst_dmem_ram_217__4_,
         mem_stage_inst_dmem_ram_217__5_, mem_stage_inst_dmem_ram_217__6_,
         mem_stage_inst_dmem_ram_217__7_, mem_stage_inst_dmem_ram_217__8_,
         mem_stage_inst_dmem_ram_217__9_, mem_stage_inst_dmem_ram_217__10_,
         mem_stage_inst_dmem_ram_217__11_, mem_stage_inst_dmem_ram_217__12_,
         mem_stage_inst_dmem_ram_217__13_, mem_stage_inst_dmem_ram_217__14_,
         mem_stage_inst_dmem_ram_217__15_, mem_stage_inst_dmem_ram_218__0_,
         mem_stage_inst_dmem_ram_218__1_, mem_stage_inst_dmem_ram_218__2_,
         mem_stage_inst_dmem_ram_218__3_, mem_stage_inst_dmem_ram_218__4_,
         mem_stage_inst_dmem_ram_218__5_, mem_stage_inst_dmem_ram_218__6_,
         mem_stage_inst_dmem_ram_218__7_, mem_stage_inst_dmem_ram_218__8_,
         mem_stage_inst_dmem_ram_218__9_, mem_stage_inst_dmem_ram_218__10_,
         mem_stage_inst_dmem_ram_218__11_, mem_stage_inst_dmem_ram_218__12_,
         mem_stage_inst_dmem_ram_218__13_, mem_stage_inst_dmem_ram_218__14_,
         mem_stage_inst_dmem_ram_218__15_, mem_stage_inst_dmem_ram_219__0_,
         mem_stage_inst_dmem_ram_219__1_, mem_stage_inst_dmem_ram_219__2_,
         mem_stage_inst_dmem_ram_219__3_, mem_stage_inst_dmem_ram_219__4_,
         mem_stage_inst_dmem_ram_219__5_, mem_stage_inst_dmem_ram_219__6_,
         mem_stage_inst_dmem_ram_219__7_, mem_stage_inst_dmem_ram_219__8_,
         mem_stage_inst_dmem_ram_219__9_, mem_stage_inst_dmem_ram_219__10_,
         mem_stage_inst_dmem_ram_219__11_, mem_stage_inst_dmem_ram_219__12_,
         mem_stage_inst_dmem_ram_219__13_, mem_stage_inst_dmem_ram_219__14_,
         mem_stage_inst_dmem_ram_219__15_, mem_stage_inst_dmem_ram_220__0_,
         mem_stage_inst_dmem_ram_220__1_, mem_stage_inst_dmem_ram_220__2_,
         mem_stage_inst_dmem_ram_220__3_, mem_stage_inst_dmem_ram_220__4_,
         mem_stage_inst_dmem_ram_220__5_, mem_stage_inst_dmem_ram_220__6_,
         mem_stage_inst_dmem_ram_220__7_, mem_stage_inst_dmem_ram_220__8_,
         mem_stage_inst_dmem_ram_220__9_, mem_stage_inst_dmem_ram_220__10_,
         mem_stage_inst_dmem_ram_220__11_, mem_stage_inst_dmem_ram_220__12_,
         mem_stage_inst_dmem_ram_220__13_, mem_stage_inst_dmem_ram_220__14_,
         mem_stage_inst_dmem_ram_220__15_, mem_stage_inst_dmem_ram_221__0_,
         mem_stage_inst_dmem_ram_221__1_, mem_stage_inst_dmem_ram_221__2_,
         mem_stage_inst_dmem_ram_221__3_, mem_stage_inst_dmem_ram_221__4_,
         mem_stage_inst_dmem_ram_221__5_, mem_stage_inst_dmem_ram_221__6_,
         mem_stage_inst_dmem_ram_221__7_, mem_stage_inst_dmem_ram_221__8_,
         mem_stage_inst_dmem_ram_221__9_, mem_stage_inst_dmem_ram_221__10_,
         mem_stage_inst_dmem_ram_221__11_, mem_stage_inst_dmem_ram_221__12_,
         mem_stage_inst_dmem_ram_221__13_, mem_stage_inst_dmem_ram_221__14_,
         mem_stage_inst_dmem_ram_221__15_, mem_stage_inst_dmem_ram_222__0_,
         mem_stage_inst_dmem_ram_222__1_, mem_stage_inst_dmem_ram_222__2_,
         mem_stage_inst_dmem_ram_222__3_, mem_stage_inst_dmem_ram_222__4_,
         mem_stage_inst_dmem_ram_222__5_, mem_stage_inst_dmem_ram_222__6_,
         mem_stage_inst_dmem_ram_222__7_, mem_stage_inst_dmem_ram_222__8_,
         mem_stage_inst_dmem_ram_222__9_, mem_stage_inst_dmem_ram_222__10_,
         mem_stage_inst_dmem_ram_222__11_, mem_stage_inst_dmem_ram_222__12_,
         mem_stage_inst_dmem_ram_222__13_, mem_stage_inst_dmem_ram_222__14_,
         mem_stage_inst_dmem_ram_222__15_, mem_stage_inst_dmem_ram_223__0_,
         mem_stage_inst_dmem_ram_223__1_, mem_stage_inst_dmem_ram_223__2_,
         mem_stage_inst_dmem_ram_223__3_, mem_stage_inst_dmem_ram_223__4_,
         mem_stage_inst_dmem_ram_223__5_, mem_stage_inst_dmem_ram_223__6_,
         mem_stage_inst_dmem_ram_223__7_, mem_stage_inst_dmem_ram_223__8_,
         mem_stage_inst_dmem_ram_223__9_, mem_stage_inst_dmem_ram_223__10_,
         mem_stage_inst_dmem_ram_223__11_, mem_stage_inst_dmem_ram_223__12_,
         mem_stage_inst_dmem_ram_223__13_, mem_stage_inst_dmem_ram_223__14_,
         mem_stage_inst_dmem_ram_223__15_, mem_stage_inst_dmem_ram_160__0_,
         mem_stage_inst_dmem_ram_160__1_, mem_stage_inst_dmem_ram_160__2_,
         mem_stage_inst_dmem_ram_160__3_, mem_stage_inst_dmem_ram_160__4_,
         mem_stage_inst_dmem_ram_160__5_, mem_stage_inst_dmem_ram_160__6_,
         mem_stage_inst_dmem_ram_160__7_, mem_stage_inst_dmem_ram_160__8_,
         mem_stage_inst_dmem_ram_160__9_, mem_stage_inst_dmem_ram_160__10_,
         mem_stage_inst_dmem_ram_160__11_, mem_stage_inst_dmem_ram_160__12_,
         mem_stage_inst_dmem_ram_160__13_, mem_stage_inst_dmem_ram_160__14_,
         mem_stage_inst_dmem_ram_160__15_, mem_stage_inst_dmem_ram_161__0_,
         mem_stage_inst_dmem_ram_161__1_, mem_stage_inst_dmem_ram_161__2_,
         mem_stage_inst_dmem_ram_161__3_, mem_stage_inst_dmem_ram_161__4_,
         mem_stage_inst_dmem_ram_161__5_, mem_stage_inst_dmem_ram_161__6_,
         mem_stage_inst_dmem_ram_161__7_, mem_stage_inst_dmem_ram_161__8_,
         mem_stage_inst_dmem_ram_161__9_, mem_stage_inst_dmem_ram_161__10_,
         mem_stage_inst_dmem_ram_161__11_, mem_stage_inst_dmem_ram_161__12_,
         mem_stage_inst_dmem_ram_161__13_, mem_stage_inst_dmem_ram_161__14_,
         mem_stage_inst_dmem_ram_161__15_, mem_stage_inst_dmem_ram_162__0_,
         mem_stage_inst_dmem_ram_162__1_, mem_stage_inst_dmem_ram_162__2_,
         mem_stage_inst_dmem_ram_162__3_, mem_stage_inst_dmem_ram_162__4_,
         mem_stage_inst_dmem_ram_162__5_, mem_stage_inst_dmem_ram_162__6_,
         mem_stage_inst_dmem_ram_162__7_, mem_stage_inst_dmem_ram_162__8_,
         mem_stage_inst_dmem_ram_162__9_, mem_stage_inst_dmem_ram_162__10_,
         mem_stage_inst_dmem_ram_162__11_, mem_stage_inst_dmem_ram_162__12_,
         mem_stage_inst_dmem_ram_162__13_, mem_stage_inst_dmem_ram_162__14_,
         mem_stage_inst_dmem_ram_162__15_, mem_stage_inst_dmem_ram_163__0_,
         mem_stage_inst_dmem_ram_163__1_, mem_stage_inst_dmem_ram_163__2_,
         mem_stage_inst_dmem_ram_163__3_, mem_stage_inst_dmem_ram_163__4_,
         mem_stage_inst_dmem_ram_163__5_, mem_stage_inst_dmem_ram_163__6_,
         mem_stage_inst_dmem_ram_163__7_, mem_stage_inst_dmem_ram_163__8_,
         mem_stage_inst_dmem_ram_163__9_, mem_stage_inst_dmem_ram_163__10_,
         mem_stage_inst_dmem_ram_163__11_, mem_stage_inst_dmem_ram_163__12_,
         mem_stage_inst_dmem_ram_163__13_, mem_stage_inst_dmem_ram_163__14_,
         mem_stage_inst_dmem_ram_163__15_, mem_stage_inst_dmem_ram_164__0_,
         mem_stage_inst_dmem_ram_164__1_, mem_stage_inst_dmem_ram_164__2_,
         mem_stage_inst_dmem_ram_164__3_, mem_stage_inst_dmem_ram_164__4_,
         mem_stage_inst_dmem_ram_164__5_, mem_stage_inst_dmem_ram_164__6_,
         mem_stage_inst_dmem_ram_164__7_, mem_stage_inst_dmem_ram_164__8_,
         mem_stage_inst_dmem_ram_164__9_, mem_stage_inst_dmem_ram_164__10_,
         mem_stage_inst_dmem_ram_164__11_, mem_stage_inst_dmem_ram_164__12_,
         mem_stage_inst_dmem_ram_164__13_, mem_stage_inst_dmem_ram_164__14_,
         mem_stage_inst_dmem_ram_164__15_, mem_stage_inst_dmem_ram_165__0_,
         mem_stage_inst_dmem_ram_165__1_, mem_stage_inst_dmem_ram_165__2_,
         mem_stage_inst_dmem_ram_165__3_, mem_stage_inst_dmem_ram_165__4_,
         mem_stage_inst_dmem_ram_165__5_, mem_stage_inst_dmem_ram_165__6_,
         mem_stage_inst_dmem_ram_165__7_, mem_stage_inst_dmem_ram_165__8_,
         mem_stage_inst_dmem_ram_165__9_, mem_stage_inst_dmem_ram_165__10_,
         mem_stage_inst_dmem_ram_165__11_, mem_stage_inst_dmem_ram_165__12_,
         mem_stage_inst_dmem_ram_165__13_, mem_stage_inst_dmem_ram_165__14_,
         mem_stage_inst_dmem_ram_165__15_, mem_stage_inst_dmem_ram_166__0_,
         mem_stage_inst_dmem_ram_166__1_, mem_stage_inst_dmem_ram_166__2_,
         mem_stage_inst_dmem_ram_166__3_, mem_stage_inst_dmem_ram_166__4_,
         mem_stage_inst_dmem_ram_166__5_, mem_stage_inst_dmem_ram_166__6_,
         mem_stage_inst_dmem_ram_166__7_, mem_stage_inst_dmem_ram_166__8_,
         mem_stage_inst_dmem_ram_166__9_, mem_stage_inst_dmem_ram_166__10_,
         mem_stage_inst_dmem_ram_166__11_, mem_stage_inst_dmem_ram_166__12_,
         mem_stage_inst_dmem_ram_166__13_, mem_stage_inst_dmem_ram_166__14_,
         mem_stage_inst_dmem_ram_166__15_, mem_stage_inst_dmem_ram_167__0_,
         mem_stage_inst_dmem_ram_167__1_, mem_stage_inst_dmem_ram_167__2_,
         mem_stage_inst_dmem_ram_167__3_, mem_stage_inst_dmem_ram_167__4_,
         mem_stage_inst_dmem_ram_167__5_, mem_stage_inst_dmem_ram_167__6_,
         mem_stage_inst_dmem_ram_167__7_, mem_stage_inst_dmem_ram_167__8_,
         mem_stage_inst_dmem_ram_167__9_, mem_stage_inst_dmem_ram_167__10_,
         mem_stage_inst_dmem_ram_167__11_, mem_stage_inst_dmem_ram_167__12_,
         mem_stage_inst_dmem_ram_167__13_, mem_stage_inst_dmem_ram_167__14_,
         mem_stage_inst_dmem_ram_167__15_, mem_stage_inst_dmem_ram_168__0_,
         mem_stage_inst_dmem_ram_168__1_, mem_stage_inst_dmem_ram_168__2_,
         mem_stage_inst_dmem_ram_168__3_, mem_stage_inst_dmem_ram_168__4_,
         mem_stage_inst_dmem_ram_168__5_, mem_stage_inst_dmem_ram_168__6_,
         mem_stage_inst_dmem_ram_168__7_, mem_stage_inst_dmem_ram_168__8_,
         mem_stage_inst_dmem_ram_168__9_, mem_stage_inst_dmem_ram_168__10_,
         mem_stage_inst_dmem_ram_168__11_, mem_stage_inst_dmem_ram_168__12_,
         mem_stage_inst_dmem_ram_168__13_, mem_stage_inst_dmem_ram_168__14_,
         mem_stage_inst_dmem_ram_168__15_, mem_stage_inst_dmem_ram_169__0_,
         mem_stage_inst_dmem_ram_169__1_, mem_stage_inst_dmem_ram_169__2_,
         mem_stage_inst_dmem_ram_169__3_, mem_stage_inst_dmem_ram_169__4_,
         mem_stage_inst_dmem_ram_169__5_, mem_stage_inst_dmem_ram_169__6_,
         mem_stage_inst_dmem_ram_169__7_, mem_stage_inst_dmem_ram_169__8_,
         mem_stage_inst_dmem_ram_169__9_, mem_stage_inst_dmem_ram_169__10_,
         mem_stage_inst_dmem_ram_169__11_, mem_stage_inst_dmem_ram_169__12_,
         mem_stage_inst_dmem_ram_169__13_, mem_stage_inst_dmem_ram_169__14_,
         mem_stage_inst_dmem_ram_169__15_, mem_stage_inst_dmem_ram_170__0_,
         mem_stage_inst_dmem_ram_170__1_, mem_stage_inst_dmem_ram_170__2_,
         mem_stage_inst_dmem_ram_170__3_, mem_stage_inst_dmem_ram_170__4_,
         mem_stage_inst_dmem_ram_170__5_, mem_stage_inst_dmem_ram_170__6_,
         mem_stage_inst_dmem_ram_170__7_, mem_stage_inst_dmem_ram_170__8_,
         mem_stage_inst_dmem_ram_170__9_, mem_stage_inst_dmem_ram_170__10_,
         mem_stage_inst_dmem_ram_170__11_, mem_stage_inst_dmem_ram_170__12_,
         mem_stage_inst_dmem_ram_170__13_, mem_stage_inst_dmem_ram_170__14_,
         mem_stage_inst_dmem_ram_170__15_, mem_stage_inst_dmem_ram_171__0_,
         mem_stage_inst_dmem_ram_171__1_, mem_stage_inst_dmem_ram_171__2_,
         mem_stage_inst_dmem_ram_171__3_, mem_stage_inst_dmem_ram_171__4_,
         mem_stage_inst_dmem_ram_171__5_, mem_stage_inst_dmem_ram_171__6_,
         mem_stage_inst_dmem_ram_171__7_, mem_stage_inst_dmem_ram_171__8_,
         mem_stage_inst_dmem_ram_171__9_, mem_stage_inst_dmem_ram_171__10_,
         mem_stage_inst_dmem_ram_171__11_, mem_stage_inst_dmem_ram_171__12_,
         mem_stage_inst_dmem_ram_171__13_, mem_stage_inst_dmem_ram_171__14_,
         mem_stage_inst_dmem_ram_171__15_, mem_stage_inst_dmem_ram_172__0_,
         mem_stage_inst_dmem_ram_172__1_, mem_stage_inst_dmem_ram_172__2_,
         mem_stage_inst_dmem_ram_172__3_, mem_stage_inst_dmem_ram_172__4_,
         mem_stage_inst_dmem_ram_172__5_, mem_stage_inst_dmem_ram_172__6_,
         mem_stage_inst_dmem_ram_172__7_, mem_stage_inst_dmem_ram_172__8_,
         mem_stage_inst_dmem_ram_172__9_, mem_stage_inst_dmem_ram_172__10_,
         mem_stage_inst_dmem_ram_172__11_, mem_stage_inst_dmem_ram_172__12_,
         mem_stage_inst_dmem_ram_172__13_, mem_stage_inst_dmem_ram_172__14_,
         mem_stage_inst_dmem_ram_172__15_, mem_stage_inst_dmem_ram_173__0_,
         mem_stage_inst_dmem_ram_173__1_, mem_stage_inst_dmem_ram_173__2_,
         mem_stage_inst_dmem_ram_173__3_, mem_stage_inst_dmem_ram_173__4_,
         mem_stage_inst_dmem_ram_173__5_, mem_stage_inst_dmem_ram_173__6_,
         mem_stage_inst_dmem_ram_173__7_, mem_stage_inst_dmem_ram_173__8_,
         mem_stage_inst_dmem_ram_173__9_, mem_stage_inst_dmem_ram_173__10_,
         mem_stage_inst_dmem_ram_173__11_, mem_stage_inst_dmem_ram_173__12_,
         mem_stage_inst_dmem_ram_173__13_, mem_stage_inst_dmem_ram_173__14_,
         mem_stage_inst_dmem_ram_173__15_, mem_stage_inst_dmem_ram_174__0_,
         mem_stage_inst_dmem_ram_174__1_, mem_stage_inst_dmem_ram_174__2_,
         mem_stage_inst_dmem_ram_174__3_, mem_stage_inst_dmem_ram_174__4_,
         mem_stage_inst_dmem_ram_174__5_, mem_stage_inst_dmem_ram_174__6_,
         mem_stage_inst_dmem_ram_174__7_, mem_stage_inst_dmem_ram_174__8_,
         mem_stage_inst_dmem_ram_174__9_, mem_stage_inst_dmem_ram_174__10_,
         mem_stage_inst_dmem_ram_174__11_, mem_stage_inst_dmem_ram_174__12_,
         mem_stage_inst_dmem_ram_174__13_, mem_stage_inst_dmem_ram_174__14_,
         mem_stage_inst_dmem_ram_174__15_, mem_stage_inst_dmem_ram_175__0_,
         mem_stage_inst_dmem_ram_175__1_, mem_stage_inst_dmem_ram_175__2_,
         mem_stage_inst_dmem_ram_175__3_, mem_stage_inst_dmem_ram_175__4_,
         mem_stage_inst_dmem_ram_175__5_, mem_stage_inst_dmem_ram_175__6_,
         mem_stage_inst_dmem_ram_175__7_, mem_stage_inst_dmem_ram_175__8_,
         mem_stage_inst_dmem_ram_175__9_, mem_stage_inst_dmem_ram_175__10_,
         mem_stage_inst_dmem_ram_175__11_, mem_stage_inst_dmem_ram_175__12_,
         mem_stage_inst_dmem_ram_175__13_, mem_stage_inst_dmem_ram_175__14_,
         mem_stage_inst_dmem_ram_175__15_, mem_stage_inst_dmem_ram_176__0_,
         mem_stage_inst_dmem_ram_176__1_, mem_stage_inst_dmem_ram_176__2_,
         mem_stage_inst_dmem_ram_176__3_, mem_stage_inst_dmem_ram_176__4_,
         mem_stage_inst_dmem_ram_176__5_, mem_stage_inst_dmem_ram_176__6_,
         mem_stage_inst_dmem_ram_176__7_, mem_stage_inst_dmem_ram_176__8_,
         mem_stage_inst_dmem_ram_176__9_, mem_stage_inst_dmem_ram_176__10_,
         mem_stage_inst_dmem_ram_176__11_, mem_stage_inst_dmem_ram_176__12_,
         mem_stage_inst_dmem_ram_176__13_, mem_stage_inst_dmem_ram_176__14_,
         mem_stage_inst_dmem_ram_176__15_, mem_stage_inst_dmem_ram_177__0_,
         mem_stage_inst_dmem_ram_177__1_, mem_stage_inst_dmem_ram_177__2_,
         mem_stage_inst_dmem_ram_177__3_, mem_stage_inst_dmem_ram_177__4_,
         mem_stage_inst_dmem_ram_177__5_, mem_stage_inst_dmem_ram_177__6_,
         mem_stage_inst_dmem_ram_177__7_, mem_stage_inst_dmem_ram_177__8_,
         mem_stage_inst_dmem_ram_177__9_, mem_stage_inst_dmem_ram_177__10_,
         mem_stage_inst_dmem_ram_177__11_, mem_stage_inst_dmem_ram_177__12_,
         mem_stage_inst_dmem_ram_177__13_, mem_stage_inst_dmem_ram_177__14_,
         mem_stage_inst_dmem_ram_177__15_, mem_stage_inst_dmem_ram_178__0_,
         mem_stage_inst_dmem_ram_178__1_, mem_stage_inst_dmem_ram_178__2_,
         mem_stage_inst_dmem_ram_178__3_, mem_stage_inst_dmem_ram_178__4_,
         mem_stage_inst_dmem_ram_178__5_, mem_stage_inst_dmem_ram_178__6_,
         mem_stage_inst_dmem_ram_178__7_, mem_stage_inst_dmem_ram_178__8_,
         mem_stage_inst_dmem_ram_178__9_, mem_stage_inst_dmem_ram_178__10_,
         mem_stage_inst_dmem_ram_178__11_, mem_stage_inst_dmem_ram_178__12_,
         mem_stage_inst_dmem_ram_178__13_, mem_stage_inst_dmem_ram_178__14_,
         mem_stage_inst_dmem_ram_178__15_, mem_stage_inst_dmem_ram_179__0_,
         mem_stage_inst_dmem_ram_179__1_, mem_stage_inst_dmem_ram_179__2_,
         mem_stage_inst_dmem_ram_179__3_, mem_stage_inst_dmem_ram_179__4_,
         mem_stage_inst_dmem_ram_179__5_, mem_stage_inst_dmem_ram_179__6_,
         mem_stage_inst_dmem_ram_179__7_, mem_stage_inst_dmem_ram_179__8_,
         mem_stage_inst_dmem_ram_179__9_, mem_stage_inst_dmem_ram_179__10_,
         mem_stage_inst_dmem_ram_179__11_, mem_stage_inst_dmem_ram_179__12_,
         mem_stage_inst_dmem_ram_179__13_, mem_stage_inst_dmem_ram_179__14_,
         mem_stage_inst_dmem_ram_179__15_, mem_stage_inst_dmem_ram_180__0_,
         mem_stage_inst_dmem_ram_180__1_, mem_stage_inst_dmem_ram_180__2_,
         mem_stage_inst_dmem_ram_180__3_, mem_stage_inst_dmem_ram_180__4_,
         mem_stage_inst_dmem_ram_180__5_, mem_stage_inst_dmem_ram_180__6_,
         mem_stage_inst_dmem_ram_180__7_, mem_stage_inst_dmem_ram_180__8_,
         mem_stage_inst_dmem_ram_180__9_, mem_stage_inst_dmem_ram_180__10_,
         mem_stage_inst_dmem_ram_180__11_, mem_stage_inst_dmem_ram_180__12_,
         mem_stage_inst_dmem_ram_180__13_, mem_stage_inst_dmem_ram_180__14_,
         mem_stage_inst_dmem_ram_180__15_, mem_stage_inst_dmem_ram_181__0_,
         mem_stage_inst_dmem_ram_181__1_, mem_stage_inst_dmem_ram_181__2_,
         mem_stage_inst_dmem_ram_181__3_, mem_stage_inst_dmem_ram_181__4_,
         mem_stage_inst_dmem_ram_181__5_, mem_stage_inst_dmem_ram_181__6_,
         mem_stage_inst_dmem_ram_181__7_, mem_stage_inst_dmem_ram_181__8_,
         mem_stage_inst_dmem_ram_181__9_, mem_stage_inst_dmem_ram_181__10_,
         mem_stage_inst_dmem_ram_181__11_, mem_stage_inst_dmem_ram_181__12_,
         mem_stage_inst_dmem_ram_181__13_, mem_stage_inst_dmem_ram_181__14_,
         mem_stage_inst_dmem_ram_181__15_, mem_stage_inst_dmem_ram_182__0_,
         mem_stage_inst_dmem_ram_182__1_, mem_stage_inst_dmem_ram_182__2_,
         mem_stage_inst_dmem_ram_182__3_, mem_stage_inst_dmem_ram_182__4_,
         mem_stage_inst_dmem_ram_182__5_, mem_stage_inst_dmem_ram_182__6_,
         mem_stage_inst_dmem_ram_182__7_, mem_stage_inst_dmem_ram_182__8_,
         mem_stage_inst_dmem_ram_182__9_, mem_stage_inst_dmem_ram_182__10_,
         mem_stage_inst_dmem_ram_182__11_, mem_stage_inst_dmem_ram_182__12_,
         mem_stage_inst_dmem_ram_182__13_, mem_stage_inst_dmem_ram_182__14_,
         mem_stage_inst_dmem_ram_182__15_, mem_stage_inst_dmem_ram_183__0_,
         mem_stage_inst_dmem_ram_183__1_, mem_stage_inst_dmem_ram_183__2_,
         mem_stage_inst_dmem_ram_183__3_, mem_stage_inst_dmem_ram_183__4_,
         mem_stage_inst_dmem_ram_183__5_, mem_stage_inst_dmem_ram_183__6_,
         mem_stage_inst_dmem_ram_183__7_, mem_stage_inst_dmem_ram_183__8_,
         mem_stage_inst_dmem_ram_183__9_, mem_stage_inst_dmem_ram_183__10_,
         mem_stage_inst_dmem_ram_183__11_, mem_stage_inst_dmem_ram_183__12_,
         mem_stage_inst_dmem_ram_183__13_, mem_stage_inst_dmem_ram_183__14_,
         mem_stage_inst_dmem_ram_183__15_, mem_stage_inst_dmem_ram_184__0_,
         mem_stage_inst_dmem_ram_184__1_, mem_stage_inst_dmem_ram_184__2_,
         mem_stage_inst_dmem_ram_184__3_, mem_stage_inst_dmem_ram_184__4_,
         mem_stage_inst_dmem_ram_184__5_, mem_stage_inst_dmem_ram_184__6_,
         mem_stage_inst_dmem_ram_184__7_, mem_stage_inst_dmem_ram_184__8_,
         mem_stage_inst_dmem_ram_184__9_, mem_stage_inst_dmem_ram_184__10_,
         mem_stage_inst_dmem_ram_184__11_, mem_stage_inst_dmem_ram_184__12_,
         mem_stage_inst_dmem_ram_184__13_, mem_stage_inst_dmem_ram_184__14_,
         mem_stage_inst_dmem_ram_184__15_, mem_stage_inst_dmem_ram_185__0_,
         mem_stage_inst_dmem_ram_185__1_, mem_stage_inst_dmem_ram_185__2_,
         mem_stage_inst_dmem_ram_185__3_, mem_stage_inst_dmem_ram_185__4_,
         mem_stage_inst_dmem_ram_185__5_, mem_stage_inst_dmem_ram_185__6_,
         mem_stage_inst_dmem_ram_185__7_, mem_stage_inst_dmem_ram_185__8_,
         mem_stage_inst_dmem_ram_185__9_, mem_stage_inst_dmem_ram_185__10_,
         mem_stage_inst_dmem_ram_185__11_, mem_stage_inst_dmem_ram_185__12_,
         mem_stage_inst_dmem_ram_185__13_, mem_stage_inst_dmem_ram_185__14_,
         mem_stage_inst_dmem_ram_185__15_, mem_stage_inst_dmem_ram_186__0_,
         mem_stage_inst_dmem_ram_186__1_, mem_stage_inst_dmem_ram_186__2_,
         mem_stage_inst_dmem_ram_186__3_, mem_stage_inst_dmem_ram_186__4_,
         mem_stage_inst_dmem_ram_186__5_, mem_stage_inst_dmem_ram_186__6_,
         mem_stage_inst_dmem_ram_186__7_, mem_stage_inst_dmem_ram_186__8_,
         mem_stage_inst_dmem_ram_186__9_, mem_stage_inst_dmem_ram_186__10_,
         mem_stage_inst_dmem_ram_186__11_, mem_stage_inst_dmem_ram_186__12_,
         mem_stage_inst_dmem_ram_186__13_, mem_stage_inst_dmem_ram_186__14_,
         mem_stage_inst_dmem_ram_186__15_, mem_stage_inst_dmem_ram_187__0_,
         mem_stage_inst_dmem_ram_187__1_, mem_stage_inst_dmem_ram_187__2_,
         mem_stage_inst_dmem_ram_187__3_, mem_stage_inst_dmem_ram_187__4_,
         mem_stage_inst_dmem_ram_187__5_, mem_stage_inst_dmem_ram_187__6_,
         mem_stage_inst_dmem_ram_187__7_, mem_stage_inst_dmem_ram_187__8_,
         mem_stage_inst_dmem_ram_187__9_, mem_stage_inst_dmem_ram_187__10_,
         mem_stage_inst_dmem_ram_187__11_, mem_stage_inst_dmem_ram_187__12_,
         mem_stage_inst_dmem_ram_187__13_, mem_stage_inst_dmem_ram_187__14_,
         mem_stage_inst_dmem_ram_187__15_, mem_stage_inst_dmem_ram_188__0_,
         mem_stage_inst_dmem_ram_188__1_, mem_stage_inst_dmem_ram_188__2_,
         mem_stage_inst_dmem_ram_188__3_, mem_stage_inst_dmem_ram_188__4_,
         mem_stage_inst_dmem_ram_188__5_, mem_stage_inst_dmem_ram_188__6_,
         mem_stage_inst_dmem_ram_188__7_, mem_stage_inst_dmem_ram_188__8_,
         mem_stage_inst_dmem_ram_188__9_, mem_stage_inst_dmem_ram_188__10_,
         mem_stage_inst_dmem_ram_188__11_, mem_stage_inst_dmem_ram_188__12_,
         mem_stage_inst_dmem_ram_188__13_, mem_stage_inst_dmem_ram_188__14_,
         mem_stage_inst_dmem_ram_188__15_, mem_stage_inst_dmem_ram_189__0_,
         mem_stage_inst_dmem_ram_189__1_, mem_stage_inst_dmem_ram_189__2_,
         mem_stage_inst_dmem_ram_189__3_, mem_stage_inst_dmem_ram_189__4_,
         mem_stage_inst_dmem_ram_189__5_, mem_stage_inst_dmem_ram_189__6_,
         mem_stage_inst_dmem_ram_189__7_, mem_stage_inst_dmem_ram_189__8_,
         mem_stage_inst_dmem_ram_189__9_, mem_stage_inst_dmem_ram_189__10_,
         mem_stage_inst_dmem_ram_189__11_, mem_stage_inst_dmem_ram_189__12_,
         mem_stage_inst_dmem_ram_189__13_, mem_stage_inst_dmem_ram_189__14_,
         mem_stage_inst_dmem_ram_189__15_, mem_stage_inst_dmem_ram_190__0_,
         mem_stage_inst_dmem_ram_190__1_, mem_stage_inst_dmem_ram_190__2_,
         mem_stage_inst_dmem_ram_190__3_, mem_stage_inst_dmem_ram_190__4_,
         mem_stage_inst_dmem_ram_190__5_, mem_stage_inst_dmem_ram_190__6_,
         mem_stage_inst_dmem_ram_190__7_, mem_stage_inst_dmem_ram_190__8_,
         mem_stage_inst_dmem_ram_190__9_, mem_stage_inst_dmem_ram_190__10_,
         mem_stage_inst_dmem_ram_190__11_, mem_stage_inst_dmem_ram_190__12_,
         mem_stage_inst_dmem_ram_190__13_, mem_stage_inst_dmem_ram_190__14_,
         mem_stage_inst_dmem_ram_190__15_, mem_stage_inst_dmem_ram_191__0_,
         mem_stage_inst_dmem_ram_191__1_, mem_stage_inst_dmem_ram_191__2_,
         mem_stage_inst_dmem_ram_191__3_, mem_stage_inst_dmem_ram_191__4_,
         mem_stage_inst_dmem_ram_191__5_, mem_stage_inst_dmem_ram_191__6_,
         mem_stage_inst_dmem_ram_191__7_, mem_stage_inst_dmem_ram_191__8_,
         mem_stage_inst_dmem_ram_191__9_, mem_stage_inst_dmem_ram_191__10_,
         mem_stage_inst_dmem_ram_191__11_, mem_stage_inst_dmem_ram_191__12_,
         mem_stage_inst_dmem_ram_191__13_, mem_stage_inst_dmem_ram_191__14_,
         mem_stage_inst_dmem_ram_191__15_, mem_stage_inst_dmem_ram_128__0_,
         mem_stage_inst_dmem_ram_128__1_, mem_stage_inst_dmem_ram_128__2_,
         mem_stage_inst_dmem_ram_128__3_, mem_stage_inst_dmem_ram_128__4_,
         mem_stage_inst_dmem_ram_128__5_, mem_stage_inst_dmem_ram_128__6_,
         mem_stage_inst_dmem_ram_128__7_, mem_stage_inst_dmem_ram_128__8_,
         mem_stage_inst_dmem_ram_128__9_, mem_stage_inst_dmem_ram_128__10_,
         mem_stage_inst_dmem_ram_128__11_, mem_stage_inst_dmem_ram_128__12_,
         mem_stage_inst_dmem_ram_128__13_, mem_stage_inst_dmem_ram_128__14_,
         mem_stage_inst_dmem_ram_128__15_, mem_stage_inst_dmem_ram_129__0_,
         mem_stage_inst_dmem_ram_129__1_, mem_stage_inst_dmem_ram_129__2_,
         mem_stage_inst_dmem_ram_129__3_, mem_stage_inst_dmem_ram_129__4_,
         mem_stage_inst_dmem_ram_129__5_, mem_stage_inst_dmem_ram_129__6_,
         mem_stage_inst_dmem_ram_129__7_, mem_stage_inst_dmem_ram_129__8_,
         mem_stage_inst_dmem_ram_129__9_, mem_stage_inst_dmem_ram_129__10_,
         mem_stage_inst_dmem_ram_129__11_, mem_stage_inst_dmem_ram_129__12_,
         mem_stage_inst_dmem_ram_129__13_, mem_stage_inst_dmem_ram_129__14_,
         mem_stage_inst_dmem_ram_129__15_, mem_stage_inst_dmem_ram_130__0_,
         mem_stage_inst_dmem_ram_130__1_, mem_stage_inst_dmem_ram_130__2_,
         mem_stage_inst_dmem_ram_130__3_, mem_stage_inst_dmem_ram_130__4_,
         mem_stage_inst_dmem_ram_130__5_, mem_stage_inst_dmem_ram_130__6_,
         mem_stage_inst_dmem_ram_130__7_, mem_stage_inst_dmem_ram_130__8_,
         mem_stage_inst_dmem_ram_130__9_, mem_stage_inst_dmem_ram_130__10_,
         mem_stage_inst_dmem_ram_130__11_, mem_stage_inst_dmem_ram_130__12_,
         mem_stage_inst_dmem_ram_130__13_, mem_stage_inst_dmem_ram_130__14_,
         mem_stage_inst_dmem_ram_130__15_, mem_stage_inst_dmem_ram_131__0_,
         mem_stage_inst_dmem_ram_131__1_, mem_stage_inst_dmem_ram_131__2_,
         mem_stage_inst_dmem_ram_131__3_, mem_stage_inst_dmem_ram_131__4_,
         mem_stage_inst_dmem_ram_131__5_, mem_stage_inst_dmem_ram_131__6_,
         mem_stage_inst_dmem_ram_131__7_, mem_stage_inst_dmem_ram_131__8_,
         mem_stage_inst_dmem_ram_131__9_, mem_stage_inst_dmem_ram_131__10_,
         mem_stage_inst_dmem_ram_131__11_, mem_stage_inst_dmem_ram_131__12_,
         mem_stage_inst_dmem_ram_131__13_, mem_stage_inst_dmem_ram_131__14_,
         mem_stage_inst_dmem_ram_131__15_, mem_stage_inst_dmem_ram_132__0_,
         mem_stage_inst_dmem_ram_132__1_, mem_stage_inst_dmem_ram_132__2_,
         mem_stage_inst_dmem_ram_132__3_, mem_stage_inst_dmem_ram_132__4_,
         mem_stage_inst_dmem_ram_132__5_, mem_stage_inst_dmem_ram_132__6_,
         mem_stage_inst_dmem_ram_132__7_, mem_stage_inst_dmem_ram_132__8_,
         mem_stage_inst_dmem_ram_132__9_, mem_stage_inst_dmem_ram_132__10_,
         mem_stage_inst_dmem_ram_132__11_, mem_stage_inst_dmem_ram_132__12_,
         mem_stage_inst_dmem_ram_132__13_, mem_stage_inst_dmem_ram_132__14_,
         mem_stage_inst_dmem_ram_132__15_, mem_stage_inst_dmem_ram_133__0_,
         mem_stage_inst_dmem_ram_133__1_, mem_stage_inst_dmem_ram_133__2_,
         mem_stage_inst_dmem_ram_133__3_, mem_stage_inst_dmem_ram_133__4_,
         mem_stage_inst_dmem_ram_133__5_, mem_stage_inst_dmem_ram_133__6_,
         mem_stage_inst_dmem_ram_133__7_, mem_stage_inst_dmem_ram_133__8_,
         mem_stage_inst_dmem_ram_133__9_, mem_stage_inst_dmem_ram_133__10_,
         mem_stage_inst_dmem_ram_133__11_, mem_stage_inst_dmem_ram_133__12_,
         mem_stage_inst_dmem_ram_133__13_, mem_stage_inst_dmem_ram_133__14_,
         mem_stage_inst_dmem_ram_133__15_, mem_stage_inst_dmem_ram_134__0_,
         mem_stage_inst_dmem_ram_134__1_, mem_stage_inst_dmem_ram_134__2_,
         mem_stage_inst_dmem_ram_134__3_, mem_stage_inst_dmem_ram_134__4_,
         mem_stage_inst_dmem_ram_134__5_, mem_stage_inst_dmem_ram_134__6_,
         mem_stage_inst_dmem_ram_134__7_, mem_stage_inst_dmem_ram_134__8_,
         mem_stage_inst_dmem_ram_134__9_, mem_stage_inst_dmem_ram_134__10_,
         mem_stage_inst_dmem_ram_134__11_, mem_stage_inst_dmem_ram_134__12_,
         mem_stage_inst_dmem_ram_134__13_, mem_stage_inst_dmem_ram_134__14_,
         mem_stage_inst_dmem_ram_134__15_, mem_stage_inst_dmem_ram_135__0_,
         mem_stage_inst_dmem_ram_135__1_, mem_stage_inst_dmem_ram_135__2_,
         mem_stage_inst_dmem_ram_135__3_, mem_stage_inst_dmem_ram_135__4_,
         mem_stage_inst_dmem_ram_135__5_, mem_stage_inst_dmem_ram_135__6_,
         mem_stage_inst_dmem_ram_135__7_, mem_stage_inst_dmem_ram_135__8_,
         mem_stage_inst_dmem_ram_135__9_, mem_stage_inst_dmem_ram_135__10_,
         mem_stage_inst_dmem_ram_135__11_, mem_stage_inst_dmem_ram_135__12_,
         mem_stage_inst_dmem_ram_135__13_, mem_stage_inst_dmem_ram_135__14_,
         mem_stage_inst_dmem_ram_135__15_, mem_stage_inst_dmem_ram_136__0_,
         mem_stage_inst_dmem_ram_136__1_, mem_stage_inst_dmem_ram_136__2_,
         mem_stage_inst_dmem_ram_136__3_, mem_stage_inst_dmem_ram_136__4_,
         mem_stage_inst_dmem_ram_136__5_, mem_stage_inst_dmem_ram_136__6_,
         mem_stage_inst_dmem_ram_136__7_, mem_stage_inst_dmem_ram_136__8_,
         mem_stage_inst_dmem_ram_136__9_, mem_stage_inst_dmem_ram_136__10_,
         mem_stage_inst_dmem_ram_136__11_, mem_stage_inst_dmem_ram_136__12_,
         mem_stage_inst_dmem_ram_136__13_, mem_stage_inst_dmem_ram_136__14_,
         mem_stage_inst_dmem_ram_136__15_, mem_stage_inst_dmem_ram_137__0_,
         mem_stage_inst_dmem_ram_137__1_, mem_stage_inst_dmem_ram_137__2_,
         mem_stage_inst_dmem_ram_137__3_, mem_stage_inst_dmem_ram_137__4_,
         mem_stage_inst_dmem_ram_137__5_, mem_stage_inst_dmem_ram_137__6_,
         mem_stage_inst_dmem_ram_137__7_, mem_stage_inst_dmem_ram_137__8_,
         mem_stage_inst_dmem_ram_137__9_, mem_stage_inst_dmem_ram_137__10_,
         mem_stage_inst_dmem_ram_137__11_, mem_stage_inst_dmem_ram_137__12_,
         mem_stage_inst_dmem_ram_137__13_, mem_stage_inst_dmem_ram_137__14_,
         mem_stage_inst_dmem_ram_137__15_, mem_stage_inst_dmem_ram_138__0_,
         mem_stage_inst_dmem_ram_138__1_, mem_stage_inst_dmem_ram_138__2_,
         mem_stage_inst_dmem_ram_138__3_, mem_stage_inst_dmem_ram_138__4_,
         mem_stage_inst_dmem_ram_138__5_, mem_stage_inst_dmem_ram_138__6_,
         mem_stage_inst_dmem_ram_138__7_, mem_stage_inst_dmem_ram_138__8_,
         mem_stage_inst_dmem_ram_138__9_, mem_stage_inst_dmem_ram_138__10_,
         mem_stage_inst_dmem_ram_138__11_, mem_stage_inst_dmem_ram_138__12_,
         mem_stage_inst_dmem_ram_138__13_, mem_stage_inst_dmem_ram_138__14_,
         mem_stage_inst_dmem_ram_138__15_, mem_stage_inst_dmem_ram_139__0_,
         mem_stage_inst_dmem_ram_139__1_, mem_stage_inst_dmem_ram_139__2_,
         mem_stage_inst_dmem_ram_139__3_, mem_stage_inst_dmem_ram_139__4_,
         mem_stage_inst_dmem_ram_139__5_, mem_stage_inst_dmem_ram_139__6_,
         mem_stage_inst_dmem_ram_139__7_, mem_stage_inst_dmem_ram_139__8_,
         mem_stage_inst_dmem_ram_139__9_, mem_stage_inst_dmem_ram_139__10_,
         mem_stage_inst_dmem_ram_139__11_, mem_stage_inst_dmem_ram_139__12_,
         mem_stage_inst_dmem_ram_139__13_, mem_stage_inst_dmem_ram_139__14_,
         mem_stage_inst_dmem_ram_139__15_, mem_stage_inst_dmem_ram_140__0_,
         mem_stage_inst_dmem_ram_140__1_, mem_stage_inst_dmem_ram_140__2_,
         mem_stage_inst_dmem_ram_140__3_, mem_stage_inst_dmem_ram_140__4_,
         mem_stage_inst_dmem_ram_140__5_, mem_stage_inst_dmem_ram_140__6_,
         mem_stage_inst_dmem_ram_140__7_, mem_stage_inst_dmem_ram_140__8_,
         mem_stage_inst_dmem_ram_140__9_, mem_stage_inst_dmem_ram_140__10_,
         mem_stage_inst_dmem_ram_140__11_, mem_stage_inst_dmem_ram_140__12_,
         mem_stage_inst_dmem_ram_140__13_, mem_stage_inst_dmem_ram_140__14_,
         mem_stage_inst_dmem_ram_140__15_, mem_stage_inst_dmem_ram_141__0_,
         mem_stage_inst_dmem_ram_141__1_, mem_stage_inst_dmem_ram_141__2_,
         mem_stage_inst_dmem_ram_141__3_, mem_stage_inst_dmem_ram_141__4_,
         mem_stage_inst_dmem_ram_141__5_, mem_stage_inst_dmem_ram_141__6_,
         mem_stage_inst_dmem_ram_141__7_, mem_stage_inst_dmem_ram_141__8_,
         mem_stage_inst_dmem_ram_141__9_, mem_stage_inst_dmem_ram_141__10_,
         mem_stage_inst_dmem_ram_141__11_, mem_stage_inst_dmem_ram_141__12_,
         mem_stage_inst_dmem_ram_141__13_, mem_stage_inst_dmem_ram_141__14_,
         mem_stage_inst_dmem_ram_141__15_, mem_stage_inst_dmem_ram_142__0_,
         mem_stage_inst_dmem_ram_142__1_, mem_stage_inst_dmem_ram_142__2_,
         mem_stage_inst_dmem_ram_142__3_, mem_stage_inst_dmem_ram_142__4_,
         mem_stage_inst_dmem_ram_142__5_, mem_stage_inst_dmem_ram_142__6_,
         mem_stage_inst_dmem_ram_142__7_, mem_stage_inst_dmem_ram_142__8_,
         mem_stage_inst_dmem_ram_142__9_, mem_stage_inst_dmem_ram_142__10_,
         mem_stage_inst_dmem_ram_142__11_, mem_stage_inst_dmem_ram_142__12_,
         mem_stage_inst_dmem_ram_142__13_, mem_stage_inst_dmem_ram_142__14_,
         mem_stage_inst_dmem_ram_142__15_, mem_stage_inst_dmem_ram_143__0_,
         mem_stage_inst_dmem_ram_143__1_, mem_stage_inst_dmem_ram_143__2_,
         mem_stage_inst_dmem_ram_143__3_, mem_stage_inst_dmem_ram_143__4_,
         mem_stage_inst_dmem_ram_143__5_, mem_stage_inst_dmem_ram_143__6_,
         mem_stage_inst_dmem_ram_143__7_, mem_stage_inst_dmem_ram_143__8_,
         mem_stage_inst_dmem_ram_143__9_, mem_stage_inst_dmem_ram_143__10_,
         mem_stage_inst_dmem_ram_143__11_, mem_stage_inst_dmem_ram_143__12_,
         mem_stage_inst_dmem_ram_143__13_, mem_stage_inst_dmem_ram_143__14_,
         mem_stage_inst_dmem_ram_143__15_, mem_stage_inst_dmem_ram_144__0_,
         mem_stage_inst_dmem_ram_144__1_, mem_stage_inst_dmem_ram_144__2_,
         mem_stage_inst_dmem_ram_144__3_, mem_stage_inst_dmem_ram_144__4_,
         mem_stage_inst_dmem_ram_144__5_, mem_stage_inst_dmem_ram_144__6_,
         mem_stage_inst_dmem_ram_144__7_, mem_stage_inst_dmem_ram_144__8_,
         mem_stage_inst_dmem_ram_144__9_, mem_stage_inst_dmem_ram_144__10_,
         mem_stage_inst_dmem_ram_144__11_, mem_stage_inst_dmem_ram_144__12_,
         mem_stage_inst_dmem_ram_144__13_, mem_stage_inst_dmem_ram_144__14_,
         mem_stage_inst_dmem_ram_144__15_, mem_stage_inst_dmem_ram_145__0_,
         mem_stage_inst_dmem_ram_145__1_, mem_stage_inst_dmem_ram_145__2_,
         mem_stage_inst_dmem_ram_145__3_, mem_stage_inst_dmem_ram_145__4_,
         mem_stage_inst_dmem_ram_145__5_, mem_stage_inst_dmem_ram_145__6_,
         mem_stage_inst_dmem_ram_145__7_, mem_stage_inst_dmem_ram_145__8_,
         mem_stage_inst_dmem_ram_145__9_, mem_stage_inst_dmem_ram_145__10_,
         mem_stage_inst_dmem_ram_145__11_, mem_stage_inst_dmem_ram_145__12_,
         mem_stage_inst_dmem_ram_145__13_, mem_stage_inst_dmem_ram_145__14_,
         mem_stage_inst_dmem_ram_145__15_, mem_stage_inst_dmem_ram_146__0_,
         mem_stage_inst_dmem_ram_146__1_, mem_stage_inst_dmem_ram_146__2_,
         mem_stage_inst_dmem_ram_146__3_, mem_stage_inst_dmem_ram_146__4_,
         mem_stage_inst_dmem_ram_146__5_, mem_stage_inst_dmem_ram_146__6_,
         mem_stage_inst_dmem_ram_146__7_, mem_stage_inst_dmem_ram_146__8_,
         mem_stage_inst_dmem_ram_146__9_, mem_stage_inst_dmem_ram_146__10_,
         mem_stage_inst_dmem_ram_146__11_, mem_stage_inst_dmem_ram_146__12_,
         mem_stage_inst_dmem_ram_146__13_, mem_stage_inst_dmem_ram_146__14_,
         mem_stage_inst_dmem_ram_146__15_, mem_stage_inst_dmem_ram_147__0_,
         mem_stage_inst_dmem_ram_147__1_, mem_stage_inst_dmem_ram_147__2_,
         mem_stage_inst_dmem_ram_147__3_, mem_stage_inst_dmem_ram_147__4_,
         mem_stage_inst_dmem_ram_147__5_, mem_stage_inst_dmem_ram_147__6_,
         mem_stage_inst_dmem_ram_147__7_, mem_stage_inst_dmem_ram_147__8_,
         mem_stage_inst_dmem_ram_147__9_, mem_stage_inst_dmem_ram_147__10_,
         mem_stage_inst_dmem_ram_147__11_, mem_stage_inst_dmem_ram_147__12_,
         mem_stage_inst_dmem_ram_147__13_, mem_stage_inst_dmem_ram_147__14_,
         mem_stage_inst_dmem_ram_147__15_, mem_stage_inst_dmem_ram_148__0_,
         mem_stage_inst_dmem_ram_148__1_, mem_stage_inst_dmem_ram_148__2_,
         mem_stage_inst_dmem_ram_148__3_, mem_stage_inst_dmem_ram_148__4_,
         mem_stage_inst_dmem_ram_148__5_, mem_stage_inst_dmem_ram_148__6_,
         mem_stage_inst_dmem_ram_148__7_, mem_stage_inst_dmem_ram_148__8_,
         mem_stage_inst_dmem_ram_148__9_, mem_stage_inst_dmem_ram_148__10_,
         mem_stage_inst_dmem_ram_148__11_, mem_stage_inst_dmem_ram_148__12_,
         mem_stage_inst_dmem_ram_148__13_, mem_stage_inst_dmem_ram_148__14_,
         mem_stage_inst_dmem_ram_148__15_, mem_stage_inst_dmem_ram_149__0_,
         mem_stage_inst_dmem_ram_149__1_, mem_stage_inst_dmem_ram_149__2_,
         mem_stage_inst_dmem_ram_149__3_, mem_stage_inst_dmem_ram_149__4_,
         mem_stage_inst_dmem_ram_149__5_, mem_stage_inst_dmem_ram_149__6_,
         mem_stage_inst_dmem_ram_149__7_, mem_stage_inst_dmem_ram_149__8_,
         mem_stage_inst_dmem_ram_149__9_, mem_stage_inst_dmem_ram_149__10_,
         mem_stage_inst_dmem_ram_149__11_, mem_stage_inst_dmem_ram_149__12_,
         mem_stage_inst_dmem_ram_149__13_, mem_stage_inst_dmem_ram_149__14_,
         mem_stage_inst_dmem_ram_149__15_, mem_stage_inst_dmem_ram_150__0_,
         mem_stage_inst_dmem_ram_150__1_, mem_stage_inst_dmem_ram_150__2_,
         mem_stage_inst_dmem_ram_150__3_, mem_stage_inst_dmem_ram_150__4_,
         mem_stage_inst_dmem_ram_150__5_, mem_stage_inst_dmem_ram_150__6_,
         mem_stage_inst_dmem_ram_150__7_, mem_stage_inst_dmem_ram_150__8_,
         mem_stage_inst_dmem_ram_150__9_, mem_stage_inst_dmem_ram_150__10_,
         mem_stage_inst_dmem_ram_150__11_, mem_stage_inst_dmem_ram_150__12_,
         mem_stage_inst_dmem_ram_150__13_, mem_stage_inst_dmem_ram_150__14_,
         mem_stage_inst_dmem_ram_150__15_, mem_stage_inst_dmem_ram_151__0_,
         mem_stage_inst_dmem_ram_151__1_, mem_stage_inst_dmem_ram_151__2_,
         mem_stage_inst_dmem_ram_151__3_, mem_stage_inst_dmem_ram_151__4_,
         mem_stage_inst_dmem_ram_151__5_, mem_stage_inst_dmem_ram_151__6_,
         mem_stage_inst_dmem_ram_151__7_, mem_stage_inst_dmem_ram_151__8_,
         mem_stage_inst_dmem_ram_151__9_, mem_stage_inst_dmem_ram_151__10_,
         mem_stage_inst_dmem_ram_151__11_, mem_stage_inst_dmem_ram_151__12_,
         mem_stage_inst_dmem_ram_151__13_, mem_stage_inst_dmem_ram_151__14_,
         mem_stage_inst_dmem_ram_151__15_, mem_stage_inst_dmem_ram_152__0_,
         mem_stage_inst_dmem_ram_152__1_, mem_stage_inst_dmem_ram_152__2_,
         mem_stage_inst_dmem_ram_152__3_, mem_stage_inst_dmem_ram_152__4_,
         mem_stage_inst_dmem_ram_152__5_, mem_stage_inst_dmem_ram_152__6_,
         mem_stage_inst_dmem_ram_152__7_, mem_stage_inst_dmem_ram_152__8_,
         mem_stage_inst_dmem_ram_152__9_, mem_stage_inst_dmem_ram_152__10_,
         mem_stage_inst_dmem_ram_152__11_, mem_stage_inst_dmem_ram_152__12_,
         mem_stage_inst_dmem_ram_152__13_, mem_stage_inst_dmem_ram_152__14_,
         mem_stage_inst_dmem_ram_152__15_, mem_stage_inst_dmem_ram_153__0_,
         mem_stage_inst_dmem_ram_153__1_, mem_stage_inst_dmem_ram_153__2_,
         mem_stage_inst_dmem_ram_153__3_, mem_stage_inst_dmem_ram_153__4_,
         mem_stage_inst_dmem_ram_153__5_, mem_stage_inst_dmem_ram_153__6_,
         mem_stage_inst_dmem_ram_153__7_, mem_stage_inst_dmem_ram_153__8_,
         mem_stage_inst_dmem_ram_153__9_, mem_stage_inst_dmem_ram_153__10_,
         mem_stage_inst_dmem_ram_153__11_, mem_stage_inst_dmem_ram_153__12_,
         mem_stage_inst_dmem_ram_153__13_, mem_stage_inst_dmem_ram_153__14_,
         mem_stage_inst_dmem_ram_153__15_, mem_stage_inst_dmem_ram_154__0_,
         mem_stage_inst_dmem_ram_154__1_, mem_stage_inst_dmem_ram_154__2_,
         mem_stage_inst_dmem_ram_154__3_, mem_stage_inst_dmem_ram_154__4_,
         mem_stage_inst_dmem_ram_154__5_, mem_stage_inst_dmem_ram_154__6_,
         mem_stage_inst_dmem_ram_154__7_, mem_stage_inst_dmem_ram_154__8_,
         mem_stage_inst_dmem_ram_154__9_, mem_stage_inst_dmem_ram_154__10_,
         mem_stage_inst_dmem_ram_154__11_, mem_stage_inst_dmem_ram_154__12_,
         mem_stage_inst_dmem_ram_154__13_, mem_stage_inst_dmem_ram_154__14_,
         mem_stage_inst_dmem_ram_154__15_, mem_stage_inst_dmem_ram_155__0_,
         mem_stage_inst_dmem_ram_155__1_, mem_stage_inst_dmem_ram_155__2_,
         mem_stage_inst_dmem_ram_155__3_, mem_stage_inst_dmem_ram_155__4_,
         mem_stage_inst_dmem_ram_155__5_, mem_stage_inst_dmem_ram_155__6_,
         mem_stage_inst_dmem_ram_155__7_, mem_stage_inst_dmem_ram_155__8_,
         mem_stage_inst_dmem_ram_155__9_, mem_stage_inst_dmem_ram_155__10_,
         mem_stage_inst_dmem_ram_155__11_, mem_stage_inst_dmem_ram_155__12_,
         mem_stage_inst_dmem_ram_155__13_, mem_stage_inst_dmem_ram_155__14_,
         mem_stage_inst_dmem_ram_155__15_, mem_stage_inst_dmem_ram_156__0_,
         mem_stage_inst_dmem_ram_156__1_, mem_stage_inst_dmem_ram_156__2_,
         mem_stage_inst_dmem_ram_156__3_, mem_stage_inst_dmem_ram_156__4_,
         mem_stage_inst_dmem_ram_156__5_, mem_stage_inst_dmem_ram_156__6_,
         mem_stage_inst_dmem_ram_156__7_, mem_stage_inst_dmem_ram_156__8_,
         mem_stage_inst_dmem_ram_156__9_, mem_stage_inst_dmem_ram_156__10_,
         mem_stage_inst_dmem_ram_156__11_, mem_stage_inst_dmem_ram_156__12_,
         mem_stage_inst_dmem_ram_156__13_, mem_stage_inst_dmem_ram_156__14_,
         mem_stage_inst_dmem_ram_156__15_, mem_stage_inst_dmem_ram_157__0_,
         mem_stage_inst_dmem_ram_157__1_, mem_stage_inst_dmem_ram_157__2_,
         mem_stage_inst_dmem_ram_157__3_, mem_stage_inst_dmem_ram_157__4_,
         mem_stage_inst_dmem_ram_157__5_, mem_stage_inst_dmem_ram_157__6_,
         mem_stage_inst_dmem_ram_157__7_, mem_stage_inst_dmem_ram_157__8_,
         mem_stage_inst_dmem_ram_157__9_, mem_stage_inst_dmem_ram_157__10_,
         mem_stage_inst_dmem_ram_157__11_, mem_stage_inst_dmem_ram_157__12_,
         mem_stage_inst_dmem_ram_157__13_, mem_stage_inst_dmem_ram_157__14_,
         mem_stage_inst_dmem_ram_157__15_, mem_stage_inst_dmem_ram_158__0_,
         mem_stage_inst_dmem_ram_158__1_, mem_stage_inst_dmem_ram_158__2_,
         mem_stage_inst_dmem_ram_158__3_, mem_stage_inst_dmem_ram_158__4_,
         mem_stage_inst_dmem_ram_158__5_, mem_stage_inst_dmem_ram_158__6_,
         mem_stage_inst_dmem_ram_158__7_, mem_stage_inst_dmem_ram_158__8_,
         mem_stage_inst_dmem_ram_158__9_, mem_stage_inst_dmem_ram_158__10_,
         mem_stage_inst_dmem_ram_158__11_, mem_stage_inst_dmem_ram_158__12_,
         mem_stage_inst_dmem_ram_158__13_, mem_stage_inst_dmem_ram_158__14_,
         mem_stage_inst_dmem_ram_158__15_, mem_stage_inst_dmem_ram_159__0_,
         mem_stage_inst_dmem_ram_159__1_, mem_stage_inst_dmem_ram_159__2_,
         mem_stage_inst_dmem_ram_159__3_, mem_stage_inst_dmem_ram_159__4_,
         mem_stage_inst_dmem_ram_159__5_, mem_stage_inst_dmem_ram_159__6_,
         mem_stage_inst_dmem_ram_159__7_, mem_stage_inst_dmem_ram_159__8_,
         mem_stage_inst_dmem_ram_159__9_, mem_stage_inst_dmem_ram_159__10_,
         mem_stage_inst_dmem_ram_159__11_, mem_stage_inst_dmem_ram_159__12_,
         mem_stage_inst_dmem_ram_159__13_, mem_stage_inst_dmem_ram_159__14_,
         mem_stage_inst_dmem_ram_159__15_, mem_stage_inst_dmem_ram_96__0_,
         mem_stage_inst_dmem_ram_96__1_, mem_stage_inst_dmem_ram_96__2_,
         mem_stage_inst_dmem_ram_96__3_, mem_stage_inst_dmem_ram_96__4_,
         mem_stage_inst_dmem_ram_96__5_, mem_stage_inst_dmem_ram_96__6_,
         mem_stage_inst_dmem_ram_96__7_, mem_stage_inst_dmem_ram_96__8_,
         mem_stage_inst_dmem_ram_96__9_, mem_stage_inst_dmem_ram_96__10_,
         mem_stage_inst_dmem_ram_96__11_, mem_stage_inst_dmem_ram_96__12_,
         mem_stage_inst_dmem_ram_96__13_, mem_stage_inst_dmem_ram_96__14_,
         mem_stage_inst_dmem_ram_96__15_, mem_stage_inst_dmem_ram_97__0_,
         mem_stage_inst_dmem_ram_97__1_, mem_stage_inst_dmem_ram_97__2_,
         mem_stage_inst_dmem_ram_97__3_, mem_stage_inst_dmem_ram_97__4_,
         mem_stage_inst_dmem_ram_97__5_, mem_stage_inst_dmem_ram_97__6_,
         mem_stage_inst_dmem_ram_97__7_, mem_stage_inst_dmem_ram_97__8_,
         mem_stage_inst_dmem_ram_97__9_, mem_stage_inst_dmem_ram_97__10_,
         mem_stage_inst_dmem_ram_97__11_, mem_stage_inst_dmem_ram_97__12_,
         mem_stage_inst_dmem_ram_97__13_, mem_stage_inst_dmem_ram_97__14_,
         mem_stage_inst_dmem_ram_97__15_, mem_stage_inst_dmem_ram_98__0_,
         mem_stage_inst_dmem_ram_98__1_, mem_stage_inst_dmem_ram_98__2_,
         mem_stage_inst_dmem_ram_98__3_, mem_stage_inst_dmem_ram_98__4_,
         mem_stage_inst_dmem_ram_98__5_, mem_stage_inst_dmem_ram_98__6_,
         mem_stage_inst_dmem_ram_98__7_, mem_stage_inst_dmem_ram_98__8_,
         mem_stage_inst_dmem_ram_98__9_, mem_stage_inst_dmem_ram_98__10_,
         mem_stage_inst_dmem_ram_98__11_, mem_stage_inst_dmem_ram_98__12_,
         mem_stage_inst_dmem_ram_98__13_, mem_stage_inst_dmem_ram_98__14_,
         mem_stage_inst_dmem_ram_98__15_, mem_stage_inst_dmem_ram_99__0_,
         mem_stage_inst_dmem_ram_99__1_, mem_stage_inst_dmem_ram_99__2_,
         mem_stage_inst_dmem_ram_99__3_, mem_stage_inst_dmem_ram_99__4_,
         mem_stage_inst_dmem_ram_99__5_, mem_stage_inst_dmem_ram_99__6_,
         mem_stage_inst_dmem_ram_99__7_, mem_stage_inst_dmem_ram_99__8_,
         mem_stage_inst_dmem_ram_99__9_, mem_stage_inst_dmem_ram_99__10_,
         mem_stage_inst_dmem_ram_99__11_, mem_stage_inst_dmem_ram_99__12_,
         mem_stage_inst_dmem_ram_99__13_, mem_stage_inst_dmem_ram_99__14_,
         mem_stage_inst_dmem_ram_99__15_, mem_stage_inst_dmem_ram_100__0_,
         mem_stage_inst_dmem_ram_100__1_, mem_stage_inst_dmem_ram_100__2_,
         mem_stage_inst_dmem_ram_100__3_, mem_stage_inst_dmem_ram_100__4_,
         mem_stage_inst_dmem_ram_100__5_, mem_stage_inst_dmem_ram_100__6_,
         mem_stage_inst_dmem_ram_100__7_, mem_stage_inst_dmem_ram_100__8_,
         mem_stage_inst_dmem_ram_100__9_, mem_stage_inst_dmem_ram_100__10_,
         mem_stage_inst_dmem_ram_100__11_, mem_stage_inst_dmem_ram_100__12_,
         mem_stage_inst_dmem_ram_100__13_, mem_stage_inst_dmem_ram_100__14_,
         mem_stage_inst_dmem_ram_100__15_, mem_stage_inst_dmem_ram_101__0_,
         mem_stage_inst_dmem_ram_101__1_, mem_stage_inst_dmem_ram_101__2_,
         mem_stage_inst_dmem_ram_101__3_, mem_stage_inst_dmem_ram_101__4_,
         mem_stage_inst_dmem_ram_101__5_, mem_stage_inst_dmem_ram_101__6_,
         mem_stage_inst_dmem_ram_101__7_, mem_stage_inst_dmem_ram_101__8_,
         mem_stage_inst_dmem_ram_101__9_, mem_stage_inst_dmem_ram_101__10_,
         mem_stage_inst_dmem_ram_101__11_, mem_stage_inst_dmem_ram_101__12_,
         mem_stage_inst_dmem_ram_101__13_, mem_stage_inst_dmem_ram_101__14_,
         mem_stage_inst_dmem_ram_101__15_, mem_stage_inst_dmem_ram_102__0_,
         mem_stage_inst_dmem_ram_102__1_, mem_stage_inst_dmem_ram_102__2_,
         mem_stage_inst_dmem_ram_102__3_, mem_stage_inst_dmem_ram_102__4_,
         mem_stage_inst_dmem_ram_102__5_, mem_stage_inst_dmem_ram_102__6_,
         mem_stage_inst_dmem_ram_102__7_, mem_stage_inst_dmem_ram_102__8_,
         mem_stage_inst_dmem_ram_102__9_, mem_stage_inst_dmem_ram_102__10_,
         mem_stage_inst_dmem_ram_102__11_, mem_stage_inst_dmem_ram_102__12_,
         mem_stage_inst_dmem_ram_102__13_, mem_stage_inst_dmem_ram_102__14_,
         mem_stage_inst_dmem_ram_102__15_, mem_stage_inst_dmem_ram_103__0_,
         mem_stage_inst_dmem_ram_103__1_, mem_stage_inst_dmem_ram_103__2_,
         mem_stage_inst_dmem_ram_103__3_, mem_stage_inst_dmem_ram_103__4_,
         mem_stage_inst_dmem_ram_103__5_, mem_stage_inst_dmem_ram_103__6_,
         mem_stage_inst_dmem_ram_103__7_, mem_stage_inst_dmem_ram_103__8_,
         mem_stage_inst_dmem_ram_103__9_, mem_stage_inst_dmem_ram_103__10_,
         mem_stage_inst_dmem_ram_103__11_, mem_stage_inst_dmem_ram_103__12_,
         mem_stage_inst_dmem_ram_103__13_, mem_stage_inst_dmem_ram_103__14_,
         mem_stage_inst_dmem_ram_103__15_, mem_stage_inst_dmem_ram_104__0_,
         mem_stage_inst_dmem_ram_104__1_, mem_stage_inst_dmem_ram_104__2_,
         mem_stage_inst_dmem_ram_104__3_, mem_stage_inst_dmem_ram_104__4_,
         mem_stage_inst_dmem_ram_104__5_, mem_stage_inst_dmem_ram_104__6_,
         mem_stage_inst_dmem_ram_104__7_, mem_stage_inst_dmem_ram_104__8_,
         mem_stage_inst_dmem_ram_104__9_, mem_stage_inst_dmem_ram_104__10_,
         mem_stage_inst_dmem_ram_104__11_, mem_stage_inst_dmem_ram_104__12_,
         mem_stage_inst_dmem_ram_104__13_, mem_stage_inst_dmem_ram_104__14_,
         mem_stage_inst_dmem_ram_104__15_, mem_stage_inst_dmem_ram_105__0_,
         mem_stage_inst_dmem_ram_105__1_, mem_stage_inst_dmem_ram_105__2_,
         mem_stage_inst_dmem_ram_105__3_, mem_stage_inst_dmem_ram_105__4_,
         mem_stage_inst_dmem_ram_105__5_, mem_stage_inst_dmem_ram_105__6_,
         mem_stage_inst_dmem_ram_105__7_, mem_stage_inst_dmem_ram_105__8_,
         mem_stage_inst_dmem_ram_105__9_, mem_stage_inst_dmem_ram_105__10_,
         mem_stage_inst_dmem_ram_105__11_, mem_stage_inst_dmem_ram_105__12_,
         mem_stage_inst_dmem_ram_105__13_, mem_stage_inst_dmem_ram_105__14_,
         mem_stage_inst_dmem_ram_105__15_, mem_stage_inst_dmem_ram_106__0_,
         mem_stage_inst_dmem_ram_106__1_, mem_stage_inst_dmem_ram_106__2_,
         mem_stage_inst_dmem_ram_106__3_, mem_stage_inst_dmem_ram_106__4_,
         mem_stage_inst_dmem_ram_106__5_, mem_stage_inst_dmem_ram_106__6_,
         mem_stage_inst_dmem_ram_106__7_, mem_stage_inst_dmem_ram_106__8_,
         mem_stage_inst_dmem_ram_106__9_, mem_stage_inst_dmem_ram_106__10_,
         mem_stage_inst_dmem_ram_106__11_, mem_stage_inst_dmem_ram_106__12_,
         mem_stage_inst_dmem_ram_106__13_, mem_stage_inst_dmem_ram_106__14_,
         mem_stage_inst_dmem_ram_106__15_, mem_stage_inst_dmem_ram_107__0_,
         mem_stage_inst_dmem_ram_107__1_, mem_stage_inst_dmem_ram_107__2_,
         mem_stage_inst_dmem_ram_107__3_, mem_stage_inst_dmem_ram_107__4_,
         mem_stage_inst_dmem_ram_107__5_, mem_stage_inst_dmem_ram_107__6_,
         mem_stage_inst_dmem_ram_107__7_, mem_stage_inst_dmem_ram_107__8_,
         mem_stage_inst_dmem_ram_107__9_, mem_stage_inst_dmem_ram_107__10_,
         mem_stage_inst_dmem_ram_107__11_, mem_stage_inst_dmem_ram_107__12_,
         mem_stage_inst_dmem_ram_107__13_, mem_stage_inst_dmem_ram_107__14_,
         mem_stage_inst_dmem_ram_107__15_, mem_stage_inst_dmem_ram_108__0_,
         mem_stage_inst_dmem_ram_108__1_, mem_stage_inst_dmem_ram_108__2_,
         mem_stage_inst_dmem_ram_108__3_, mem_stage_inst_dmem_ram_108__4_,
         mem_stage_inst_dmem_ram_108__5_, mem_stage_inst_dmem_ram_108__6_,
         mem_stage_inst_dmem_ram_108__7_, mem_stage_inst_dmem_ram_108__8_,
         mem_stage_inst_dmem_ram_108__9_, mem_stage_inst_dmem_ram_108__10_,
         mem_stage_inst_dmem_ram_108__11_, mem_stage_inst_dmem_ram_108__12_,
         mem_stage_inst_dmem_ram_108__13_, mem_stage_inst_dmem_ram_108__14_,
         mem_stage_inst_dmem_ram_108__15_, mem_stage_inst_dmem_ram_109__0_,
         mem_stage_inst_dmem_ram_109__1_, mem_stage_inst_dmem_ram_109__2_,
         mem_stage_inst_dmem_ram_109__3_, mem_stage_inst_dmem_ram_109__4_,
         mem_stage_inst_dmem_ram_109__5_, mem_stage_inst_dmem_ram_109__6_,
         mem_stage_inst_dmem_ram_109__7_, mem_stage_inst_dmem_ram_109__8_,
         mem_stage_inst_dmem_ram_109__9_, mem_stage_inst_dmem_ram_109__10_,
         mem_stage_inst_dmem_ram_109__11_, mem_stage_inst_dmem_ram_109__12_,
         mem_stage_inst_dmem_ram_109__13_, mem_stage_inst_dmem_ram_109__14_,
         mem_stage_inst_dmem_ram_109__15_, mem_stage_inst_dmem_ram_110__0_,
         mem_stage_inst_dmem_ram_110__1_, mem_stage_inst_dmem_ram_110__2_,
         mem_stage_inst_dmem_ram_110__3_, mem_stage_inst_dmem_ram_110__4_,
         mem_stage_inst_dmem_ram_110__5_, mem_stage_inst_dmem_ram_110__6_,
         mem_stage_inst_dmem_ram_110__7_, mem_stage_inst_dmem_ram_110__8_,
         mem_stage_inst_dmem_ram_110__9_, mem_stage_inst_dmem_ram_110__10_,
         mem_stage_inst_dmem_ram_110__11_, mem_stage_inst_dmem_ram_110__12_,
         mem_stage_inst_dmem_ram_110__13_, mem_stage_inst_dmem_ram_110__14_,
         mem_stage_inst_dmem_ram_110__15_, mem_stage_inst_dmem_ram_111__0_,
         mem_stage_inst_dmem_ram_111__1_, mem_stage_inst_dmem_ram_111__2_,
         mem_stage_inst_dmem_ram_111__3_, mem_stage_inst_dmem_ram_111__4_,
         mem_stage_inst_dmem_ram_111__5_, mem_stage_inst_dmem_ram_111__6_,
         mem_stage_inst_dmem_ram_111__7_, mem_stage_inst_dmem_ram_111__8_,
         mem_stage_inst_dmem_ram_111__9_, mem_stage_inst_dmem_ram_111__10_,
         mem_stage_inst_dmem_ram_111__11_, mem_stage_inst_dmem_ram_111__12_,
         mem_stage_inst_dmem_ram_111__13_, mem_stage_inst_dmem_ram_111__14_,
         mem_stage_inst_dmem_ram_111__15_, mem_stage_inst_dmem_ram_112__0_,
         mem_stage_inst_dmem_ram_112__1_, mem_stage_inst_dmem_ram_112__2_,
         mem_stage_inst_dmem_ram_112__3_, mem_stage_inst_dmem_ram_112__4_,
         mem_stage_inst_dmem_ram_112__5_, mem_stage_inst_dmem_ram_112__6_,
         mem_stage_inst_dmem_ram_112__7_, mem_stage_inst_dmem_ram_112__8_,
         mem_stage_inst_dmem_ram_112__9_, mem_stage_inst_dmem_ram_112__10_,
         mem_stage_inst_dmem_ram_112__11_, mem_stage_inst_dmem_ram_112__12_,
         mem_stage_inst_dmem_ram_112__13_, mem_stage_inst_dmem_ram_112__14_,
         mem_stage_inst_dmem_ram_112__15_, mem_stage_inst_dmem_ram_113__0_,
         mem_stage_inst_dmem_ram_113__1_, mem_stage_inst_dmem_ram_113__2_,
         mem_stage_inst_dmem_ram_113__3_, mem_stage_inst_dmem_ram_113__4_,
         mem_stage_inst_dmem_ram_113__5_, mem_stage_inst_dmem_ram_113__6_,
         mem_stage_inst_dmem_ram_113__7_, mem_stage_inst_dmem_ram_113__8_,
         mem_stage_inst_dmem_ram_113__9_, mem_stage_inst_dmem_ram_113__10_,
         mem_stage_inst_dmem_ram_113__11_, mem_stage_inst_dmem_ram_113__12_,
         mem_stage_inst_dmem_ram_113__13_, mem_stage_inst_dmem_ram_113__14_,
         mem_stage_inst_dmem_ram_113__15_, mem_stage_inst_dmem_ram_114__0_,
         mem_stage_inst_dmem_ram_114__1_, mem_stage_inst_dmem_ram_114__2_,
         mem_stage_inst_dmem_ram_114__3_, mem_stage_inst_dmem_ram_114__4_,
         mem_stage_inst_dmem_ram_114__5_, mem_stage_inst_dmem_ram_114__6_,
         mem_stage_inst_dmem_ram_114__7_, mem_stage_inst_dmem_ram_114__8_,
         mem_stage_inst_dmem_ram_114__9_, mem_stage_inst_dmem_ram_114__10_,
         mem_stage_inst_dmem_ram_114__11_, mem_stage_inst_dmem_ram_114__12_,
         mem_stage_inst_dmem_ram_114__13_, mem_stage_inst_dmem_ram_114__14_,
         mem_stage_inst_dmem_ram_114__15_, mem_stage_inst_dmem_ram_115__0_,
         mem_stage_inst_dmem_ram_115__1_, mem_stage_inst_dmem_ram_115__2_,
         mem_stage_inst_dmem_ram_115__3_, mem_stage_inst_dmem_ram_115__4_,
         mem_stage_inst_dmem_ram_115__5_, mem_stage_inst_dmem_ram_115__6_,
         mem_stage_inst_dmem_ram_115__7_, mem_stage_inst_dmem_ram_115__8_,
         mem_stage_inst_dmem_ram_115__9_, mem_stage_inst_dmem_ram_115__10_,
         mem_stage_inst_dmem_ram_115__11_, mem_stage_inst_dmem_ram_115__12_,
         mem_stage_inst_dmem_ram_115__13_, mem_stage_inst_dmem_ram_115__14_,
         mem_stage_inst_dmem_ram_115__15_, mem_stage_inst_dmem_ram_116__0_,
         mem_stage_inst_dmem_ram_116__1_, mem_stage_inst_dmem_ram_116__2_,
         mem_stage_inst_dmem_ram_116__3_, mem_stage_inst_dmem_ram_116__4_,
         mem_stage_inst_dmem_ram_116__5_, mem_stage_inst_dmem_ram_116__6_,
         mem_stage_inst_dmem_ram_116__7_, mem_stage_inst_dmem_ram_116__8_,
         mem_stage_inst_dmem_ram_116__9_, mem_stage_inst_dmem_ram_116__10_,
         mem_stage_inst_dmem_ram_116__11_, mem_stage_inst_dmem_ram_116__12_,
         mem_stage_inst_dmem_ram_116__13_, mem_stage_inst_dmem_ram_116__14_,
         mem_stage_inst_dmem_ram_116__15_, mem_stage_inst_dmem_ram_117__0_,
         mem_stage_inst_dmem_ram_117__1_, mem_stage_inst_dmem_ram_117__2_,
         mem_stage_inst_dmem_ram_117__3_, mem_stage_inst_dmem_ram_117__4_,
         mem_stage_inst_dmem_ram_117__5_, mem_stage_inst_dmem_ram_117__6_,
         mem_stage_inst_dmem_ram_117__7_, mem_stage_inst_dmem_ram_117__8_,
         mem_stage_inst_dmem_ram_117__9_, mem_stage_inst_dmem_ram_117__10_,
         mem_stage_inst_dmem_ram_117__11_, mem_stage_inst_dmem_ram_117__12_,
         mem_stage_inst_dmem_ram_117__13_, mem_stage_inst_dmem_ram_117__14_,
         mem_stage_inst_dmem_ram_117__15_, mem_stage_inst_dmem_ram_118__0_,
         mem_stage_inst_dmem_ram_118__1_, mem_stage_inst_dmem_ram_118__2_,
         mem_stage_inst_dmem_ram_118__3_, mem_stage_inst_dmem_ram_118__4_,
         mem_stage_inst_dmem_ram_118__5_, mem_stage_inst_dmem_ram_118__6_,
         mem_stage_inst_dmem_ram_118__7_, mem_stage_inst_dmem_ram_118__8_,
         mem_stage_inst_dmem_ram_118__9_, mem_stage_inst_dmem_ram_118__10_,
         mem_stage_inst_dmem_ram_118__11_, mem_stage_inst_dmem_ram_118__12_,
         mem_stage_inst_dmem_ram_118__13_, mem_stage_inst_dmem_ram_118__14_,
         mem_stage_inst_dmem_ram_118__15_, mem_stage_inst_dmem_ram_119__0_,
         mem_stage_inst_dmem_ram_119__1_, mem_stage_inst_dmem_ram_119__2_,
         mem_stage_inst_dmem_ram_119__3_, mem_stage_inst_dmem_ram_119__4_,
         mem_stage_inst_dmem_ram_119__5_, mem_stage_inst_dmem_ram_119__6_,
         mem_stage_inst_dmem_ram_119__7_, mem_stage_inst_dmem_ram_119__8_,
         mem_stage_inst_dmem_ram_119__9_, mem_stage_inst_dmem_ram_119__10_,
         mem_stage_inst_dmem_ram_119__11_, mem_stage_inst_dmem_ram_119__12_,
         mem_stage_inst_dmem_ram_119__13_, mem_stage_inst_dmem_ram_119__14_,
         mem_stage_inst_dmem_ram_119__15_, mem_stage_inst_dmem_ram_120__0_,
         mem_stage_inst_dmem_ram_120__1_, mem_stage_inst_dmem_ram_120__2_,
         mem_stage_inst_dmem_ram_120__3_, mem_stage_inst_dmem_ram_120__4_,
         mem_stage_inst_dmem_ram_120__5_, mem_stage_inst_dmem_ram_120__6_,
         mem_stage_inst_dmem_ram_120__7_, mem_stage_inst_dmem_ram_120__8_,
         mem_stage_inst_dmem_ram_120__9_, mem_stage_inst_dmem_ram_120__10_,
         mem_stage_inst_dmem_ram_120__11_, mem_stage_inst_dmem_ram_120__12_,
         mem_stage_inst_dmem_ram_120__13_, mem_stage_inst_dmem_ram_120__14_,
         mem_stage_inst_dmem_ram_120__15_, mem_stage_inst_dmem_ram_121__0_,
         mem_stage_inst_dmem_ram_121__1_, mem_stage_inst_dmem_ram_121__2_,
         mem_stage_inst_dmem_ram_121__3_, mem_stage_inst_dmem_ram_121__4_,
         mem_stage_inst_dmem_ram_121__5_, mem_stage_inst_dmem_ram_121__6_,
         mem_stage_inst_dmem_ram_121__7_, mem_stage_inst_dmem_ram_121__8_,
         mem_stage_inst_dmem_ram_121__9_, mem_stage_inst_dmem_ram_121__10_,
         mem_stage_inst_dmem_ram_121__11_, mem_stage_inst_dmem_ram_121__12_,
         mem_stage_inst_dmem_ram_121__13_, mem_stage_inst_dmem_ram_121__14_,
         mem_stage_inst_dmem_ram_121__15_, mem_stage_inst_dmem_ram_122__0_,
         mem_stage_inst_dmem_ram_122__1_, mem_stage_inst_dmem_ram_122__2_,
         mem_stage_inst_dmem_ram_122__3_, mem_stage_inst_dmem_ram_122__4_,
         mem_stage_inst_dmem_ram_122__5_, mem_stage_inst_dmem_ram_122__6_,
         mem_stage_inst_dmem_ram_122__7_, mem_stage_inst_dmem_ram_122__8_,
         mem_stage_inst_dmem_ram_122__9_, mem_stage_inst_dmem_ram_122__10_,
         mem_stage_inst_dmem_ram_122__11_, mem_stage_inst_dmem_ram_122__12_,
         mem_stage_inst_dmem_ram_122__13_, mem_stage_inst_dmem_ram_122__14_,
         mem_stage_inst_dmem_ram_122__15_, mem_stage_inst_dmem_ram_123__0_,
         mem_stage_inst_dmem_ram_123__1_, mem_stage_inst_dmem_ram_123__2_,
         mem_stage_inst_dmem_ram_123__3_, mem_stage_inst_dmem_ram_123__4_,
         mem_stage_inst_dmem_ram_123__5_, mem_stage_inst_dmem_ram_123__6_,
         mem_stage_inst_dmem_ram_123__7_, mem_stage_inst_dmem_ram_123__8_,
         mem_stage_inst_dmem_ram_123__9_, mem_stage_inst_dmem_ram_123__10_,
         mem_stage_inst_dmem_ram_123__11_, mem_stage_inst_dmem_ram_123__12_,
         mem_stage_inst_dmem_ram_123__13_, mem_stage_inst_dmem_ram_123__14_,
         mem_stage_inst_dmem_ram_123__15_, mem_stage_inst_dmem_ram_124__0_,
         mem_stage_inst_dmem_ram_124__1_, mem_stage_inst_dmem_ram_124__2_,
         mem_stage_inst_dmem_ram_124__3_, mem_stage_inst_dmem_ram_124__4_,
         mem_stage_inst_dmem_ram_124__5_, mem_stage_inst_dmem_ram_124__6_,
         mem_stage_inst_dmem_ram_124__7_, mem_stage_inst_dmem_ram_124__8_,
         mem_stage_inst_dmem_ram_124__9_, mem_stage_inst_dmem_ram_124__10_,
         mem_stage_inst_dmem_ram_124__11_, mem_stage_inst_dmem_ram_124__12_,
         mem_stage_inst_dmem_ram_124__13_, mem_stage_inst_dmem_ram_124__14_,
         mem_stage_inst_dmem_ram_124__15_, mem_stage_inst_dmem_ram_125__0_,
         mem_stage_inst_dmem_ram_125__1_, mem_stage_inst_dmem_ram_125__2_,
         mem_stage_inst_dmem_ram_125__3_, mem_stage_inst_dmem_ram_125__4_,
         mem_stage_inst_dmem_ram_125__5_, mem_stage_inst_dmem_ram_125__6_,
         mem_stage_inst_dmem_ram_125__7_, mem_stage_inst_dmem_ram_125__8_,
         mem_stage_inst_dmem_ram_125__9_, mem_stage_inst_dmem_ram_125__10_,
         mem_stage_inst_dmem_ram_125__11_, mem_stage_inst_dmem_ram_125__12_,
         mem_stage_inst_dmem_ram_125__13_, mem_stage_inst_dmem_ram_125__14_,
         mem_stage_inst_dmem_ram_125__15_, mem_stage_inst_dmem_ram_126__0_,
         mem_stage_inst_dmem_ram_126__1_, mem_stage_inst_dmem_ram_126__2_,
         mem_stage_inst_dmem_ram_126__3_, mem_stage_inst_dmem_ram_126__4_,
         mem_stage_inst_dmem_ram_126__5_, mem_stage_inst_dmem_ram_126__6_,
         mem_stage_inst_dmem_ram_126__7_, mem_stage_inst_dmem_ram_126__8_,
         mem_stage_inst_dmem_ram_126__9_, mem_stage_inst_dmem_ram_126__10_,
         mem_stage_inst_dmem_ram_126__11_, mem_stage_inst_dmem_ram_126__12_,
         mem_stage_inst_dmem_ram_126__13_, mem_stage_inst_dmem_ram_126__14_,
         mem_stage_inst_dmem_ram_126__15_, mem_stage_inst_dmem_ram_127__0_,
         mem_stage_inst_dmem_ram_127__1_, mem_stage_inst_dmem_ram_127__2_,
         mem_stage_inst_dmem_ram_127__3_, mem_stage_inst_dmem_ram_127__4_,
         mem_stage_inst_dmem_ram_127__5_, mem_stage_inst_dmem_ram_127__6_,
         mem_stage_inst_dmem_ram_127__7_, mem_stage_inst_dmem_ram_127__8_,
         mem_stage_inst_dmem_ram_127__9_, mem_stage_inst_dmem_ram_127__10_,
         mem_stage_inst_dmem_ram_127__11_, mem_stage_inst_dmem_ram_127__12_,
         mem_stage_inst_dmem_ram_127__13_, mem_stage_inst_dmem_ram_127__14_,
         mem_stage_inst_dmem_ram_127__15_, mem_stage_inst_dmem_ram_64__0_,
         mem_stage_inst_dmem_ram_64__1_, mem_stage_inst_dmem_ram_64__2_,
         mem_stage_inst_dmem_ram_64__3_, mem_stage_inst_dmem_ram_64__4_,
         mem_stage_inst_dmem_ram_64__5_, mem_stage_inst_dmem_ram_64__6_,
         mem_stage_inst_dmem_ram_64__7_, mem_stage_inst_dmem_ram_64__8_,
         mem_stage_inst_dmem_ram_64__9_, mem_stage_inst_dmem_ram_64__10_,
         mem_stage_inst_dmem_ram_64__11_, mem_stage_inst_dmem_ram_64__12_,
         mem_stage_inst_dmem_ram_64__13_, mem_stage_inst_dmem_ram_64__14_,
         mem_stage_inst_dmem_ram_64__15_, mem_stage_inst_dmem_ram_65__0_,
         mem_stage_inst_dmem_ram_65__1_, mem_stage_inst_dmem_ram_65__2_,
         mem_stage_inst_dmem_ram_65__3_, mem_stage_inst_dmem_ram_65__4_,
         mem_stage_inst_dmem_ram_65__5_, mem_stage_inst_dmem_ram_65__6_,
         mem_stage_inst_dmem_ram_65__7_, mem_stage_inst_dmem_ram_65__8_,
         mem_stage_inst_dmem_ram_65__9_, mem_stage_inst_dmem_ram_65__10_,
         mem_stage_inst_dmem_ram_65__11_, mem_stage_inst_dmem_ram_65__12_,
         mem_stage_inst_dmem_ram_65__13_, mem_stage_inst_dmem_ram_65__14_,
         mem_stage_inst_dmem_ram_65__15_, mem_stage_inst_dmem_ram_66__0_,
         mem_stage_inst_dmem_ram_66__1_, mem_stage_inst_dmem_ram_66__2_,
         mem_stage_inst_dmem_ram_66__3_, mem_stage_inst_dmem_ram_66__4_,
         mem_stage_inst_dmem_ram_66__5_, mem_stage_inst_dmem_ram_66__6_,
         mem_stage_inst_dmem_ram_66__7_, mem_stage_inst_dmem_ram_66__8_,
         mem_stage_inst_dmem_ram_66__9_, mem_stage_inst_dmem_ram_66__10_,
         mem_stage_inst_dmem_ram_66__11_, mem_stage_inst_dmem_ram_66__12_,
         mem_stage_inst_dmem_ram_66__13_, mem_stage_inst_dmem_ram_66__14_,
         mem_stage_inst_dmem_ram_66__15_, mem_stage_inst_dmem_ram_67__0_,
         mem_stage_inst_dmem_ram_67__1_, mem_stage_inst_dmem_ram_67__2_,
         mem_stage_inst_dmem_ram_67__3_, mem_stage_inst_dmem_ram_67__4_,
         mem_stage_inst_dmem_ram_67__5_, mem_stage_inst_dmem_ram_67__6_,
         mem_stage_inst_dmem_ram_67__7_, mem_stage_inst_dmem_ram_67__8_,
         mem_stage_inst_dmem_ram_67__9_, mem_stage_inst_dmem_ram_67__10_,
         mem_stage_inst_dmem_ram_67__11_, mem_stage_inst_dmem_ram_67__12_,
         mem_stage_inst_dmem_ram_67__13_, mem_stage_inst_dmem_ram_67__14_,
         mem_stage_inst_dmem_ram_67__15_, mem_stage_inst_dmem_ram_68__0_,
         mem_stage_inst_dmem_ram_68__1_, mem_stage_inst_dmem_ram_68__2_,
         mem_stage_inst_dmem_ram_68__3_, mem_stage_inst_dmem_ram_68__4_,
         mem_stage_inst_dmem_ram_68__5_, mem_stage_inst_dmem_ram_68__6_,
         mem_stage_inst_dmem_ram_68__7_, mem_stage_inst_dmem_ram_68__8_,
         mem_stage_inst_dmem_ram_68__9_, mem_stage_inst_dmem_ram_68__10_,
         mem_stage_inst_dmem_ram_68__11_, mem_stage_inst_dmem_ram_68__12_,
         mem_stage_inst_dmem_ram_68__13_, mem_stage_inst_dmem_ram_68__14_,
         mem_stage_inst_dmem_ram_68__15_, mem_stage_inst_dmem_ram_69__0_,
         mem_stage_inst_dmem_ram_69__1_, mem_stage_inst_dmem_ram_69__2_,
         mem_stage_inst_dmem_ram_69__3_, mem_stage_inst_dmem_ram_69__4_,
         mem_stage_inst_dmem_ram_69__5_, mem_stage_inst_dmem_ram_69__6_,
         mem_stage_inst_dmem_ram_69__7_, mem_stage_inst_dmem_ram_69__8_,
         mem_stage_inst_dmem_ram_69__9_, mem_stage_inst_dmem_ram_69__10_,
         mem_stage_inst_dmem_ram_69__11_, mem_stage_inst_dmem_ram_69__12_,
         mem_stage_inst_dmem_ram_69__13_, mem_stage_inst_dmem_ram_69__14_,
         mem_stage_inst_dmem_ram_69__15_, mem_stage_inst_dmem_ram_70__0_,
         mem_stage_inst_dmem_ram_70__1_, mem_stage_inst_dmem_ram_70__2_,
         mem_stage_inst_dmem_ram_70__3_, mem_stage_inst_dmem_ram_70__4_,
         mem_stage_inst_dmem_ram_70__5_, mem_stage_inst_dmem_ram_70__6_,
         mem_stage_inst_dmem_ram_70__7_, mem_stage_inst_dmem_ram_70__8_,
         mem_stage_inst_dmem_ram_70__9_, mem_stage_inst_dmem_ram_70__10_,
         mem_stage_inst_dmem_ram_70__11_, mem_stage_inst_dmem_ram_70__12_,
         mem_stage_inst_dmem_ram_70__13_, mem_stage_inst_dmem_ram_70__14_,
         mem_stage_inst_dmem_ram_70__15_, mem_stage_inst_dmem_ram_71__0_,
         mem_stage_inst_dmem_ram_71__1_, mem_stage_inst_dmem_ram_71__2_,
         mem_stage_inst_dmem_ram_71__3_, mem_stage_inst_dmem_ram_71__4_,
         mem_stage_inst_dmem_ram_71__5_, mem_stage_inst_dmem_ram_71__6_,
         mem_stage_inst_dmem_ram_71__7_, mem_stage_inst_dmem_ram_71__8_,
         mem_stage_inst_dmem_ram_71__9_, mem_stage_inst_dmem_ram_71__10_,
         mem_stage_inst_dmem_ram_71__11_, mem_stage_inst_dmem_ram_71__12_,
         mem_stage_inst_dmem_ram_71__13_, mem_stage_inst_dmem_ram_71__14_,
         mem_stage_inst_dmem_ram_71__15_, mem_stage_inst_dmem_ram_72__0_,
         mem_stage_inst_dmem_ram_72__1_, mem_stage_inst_dmem_ram_72__2_,
         mem_stage_inst_dmem_ram_72__3_, mem_stage_inst_dmem_ram_72__4_,
         mem_stage_inst_dmem_ram_72__5_, mem_stage_inst_dmem_ram_72__6_,
         mem_stage_inst_dmem_ram_72__7_, mem_stage_inst_dmem_ram_72__8_,
         mem_stage_inst_dmem_ram_72__9_, mem_stage_inst_dmem_ram_72__10_,
         mem_stage_inst_dmem_ram_72__11_, mem_stage_inst_dmem_ram_72__12_,
         mem_stage_inst_dmem_ram_72__13_, mem_stage_inst_dmem_ram_72__14_,
         mem_stage_inst_dmem_ram_72__15_, mem_stage_inst_dmem_ram_73__0_,
         mem_stage_inst_dmem_ram_73__1_, mem_stage_inst_dmem_ram_73__2_,
         mem_stage_inst_dmem_ram_73__3_, mem_stage_inst_dmem_ram_73__4_,
         mem_stage_inst_dmem_ram_73__5_, mem_stage_inst_dmem_ram_73__6_,
         mem_stage_inst_dmem_ram_73__7_, mem_stage_inst_dmem_ram_73__8_,
         mem_stage_inst_dmem_ram_73__9_, mem_stage_inst_dmem_ram_73__10_,
         mem_stage_inst_dmem_ram_73__11_, mem_stage_inst_dmem_ram_73__12_,
         mem_stage_inst_dmem_ram_73__13_, mem_stage_inst_dmem_ram_73__14_,
         mem_stage_inst_dmem_ram_73__15_, mem_stage_inst_dmem_ram_74__0_,
         mem_stage_inst_dmem_ram_74__1_, mem_stage_inst_dmem_ram_74__2_,
         mem_stage_inst_dmem_ram_74__3_, mem_stage_inst_dmem_ram_74__4_,
         mem_stage_inst_dmem_ram_74__5_, mem_stage_inst_dmem_ram_74__6_,
         mem_stage_inst_dmem_ram_74__7_, mem_stage_inst_dmem_ram_74__8_,
         mem_stage_inst_dmem_ram_74__9_, mem_stage_inst_dmem_ram_74__10_,
         mem_stage_inst_dmem_ram_74__11_, mem_stage_inst_dmem_ram_74__12_,
         mem_stage_inst_dmem_ram_74__13_, mem_stage_inst_dmem_ram_74__14_,
         mem_stage_inst_dmem_ram_74__15_, mem_stage_inst_dmem_ram_75__0_,
         mem_stage_inst_dmem_ram_75__1_, mem_stage_inst_dmem_ram_75__2_,
         mem_stage_inst_dmem_ram_75__3_, mem_stage_inst_dmem_ram_75__4_,
         mem_stage_inst_dmem_ram_75__5_, mem_stage_inst_dmem_ram_75__6_,
         mem_stage_inst_dmem_ram_75__7_, mem_stage_inst_dmem_ram_75__8_,
         mem_stage_inst_dmem_ram_75__9_, mem_stage_inst_dmem_ram_75__10_,
         mem_stage_inst_dmem_ram_75__11_, mem_stage_inst_dmem_ram_75__12_,
         mem_stage_inst_dmem_ram_75__13_, mem_stage_inst_dmem_ram_75__14_,
         mem_stage_inst_dmem_ram_75__15_, mem_stage_inst_dmem_ram_76__0_,
         mem_stage_inst_dmem_ram_76__1_, mem_stage_inst_dmem_ram_76__2_,
         mem_stage_inst_dmem_ram_76__3_, mem_stage_inst_dmem_ram_76__4_,
         mem_stage_inst_dmem_ram_76__5_, mem_stage_inst_dmem_ram_76__6_,
         mem_stage_inst_dmem_ram_76__7_, mem_stage_inst_dmem_ram_76__8_,
         mem_stage_inst_dmem_ram_76__9_, mem_stage_inst_dmem_ram_76__10_,
         mem_stage_inst_dmem_ram_76__11_, mem_stage_inst_dmem_ram_76__12_,
         mem_stage_inst_dmem_ram_76__13_, mem_stage_inst_dmem_ram_76__14_,
         mem_stage_inst_dmem_ram_76__15_, mem_stage_inst_dmem_ram_77__0_,
         mem_stage_inst_dmem_ram_77__1_, mem_stage_inst_dmem_ram_77__2_,
         mem_stage_inst_dmem_ram_77__3_, mem_stage_inst_dmem_ram_77__4_,
         mem_stage_inst_dmem_ram_77__5_, mem_stage_inst_dmem_ram_77__6_,
         mem_stage_inst_dmem_ram_77__7_, mem_stage_inst_dmem_ram_77__8_,
         mem_stage_inst_dmem_ram_77__9_, mem_stage_inst_dmem_ram_77__10_,
         mem_stage_inst_dmem_ram_77__11_, mem_stage_inst_dmem_ram_77__12_,
         mem_stage_inst_dmem_ram_77__13_, mem_stage_inst_dmem_ram_77__14_,
         mem_stage_inst_dmem_ram_77__15_, mem_stage_inst_dmem_ram_78__0_,
         mem_stage_inst_dmem_ram_78__1_, mem_stage_inst_dmem_ram_78__2_,
         mem_stage_inst_dmem_ram_78__3_, mem_stage_inst_dmem_ram_78__4_,
         mem_stage_inst_dmem_ram_78__5_, mem_stage_inst_dmem_ram_78__6_,
         mem_stage_inst_dmem_ram_78__7_, mem_stage_inst_dmem_ram_78__8_,
         mem_stage_inst_dmem_ram_78__9_, mem_stage_inst_dmem_ram_78__10_,
         mem_stage_inst_dmem_ram_78__11_, mem_stage_inst_dmem_ram_78__12_,
         mem_stage_inst_dmem_ram_78__13_, mem_stage_inst_dmem_ram_78__14_,
         mem_stage_inst_dmem_ram_78__15_, mem_stage_inst_dmem_ram_79__0_,
         mem_stage_inst_dmem_ram_79__1_, mem_stage_inst_dmem_ram_79__2_,
         mem_stage_inst_dmem_ram_79__3_, mem_stage_inst_dmem_ram_79__4_,
         mem_stage_inst_dmem_ram_79__5_, mem_stage_inst_dmem_ram_79__6_,
         mem_stage_inst_dmem_ram_79__7_, mem_stage_inst_dmem_ram_79__8_,
         mem_stage_inst_dmem_ram_79__9_, mem_stage_inst_dmem_ram_79__10_,
         mem_stage_inst_dmem_ram_79__11_, mem_stage_inst_dmem_ram_79__12_,
         mem_stage_inst_dmem_ram_79__13_, mem_stage_inst_dmem_ram_79__14_,
         mem_stage_inst_dmem_ram_79__15_, mem_stage_inst_dmem_ram_80__0_,
         mem_stage_inst_dmem_ram_80__1_, mem_stage_inst_dmem_ram_80__2_,
         mem_stage_inst_dmem_ram_80__3_, mem_stage_inst_dmem_ram_80__4_,
         mem_stage_inst_dmem_ram_80__5_, mem_stage_inst_dmem_ram_80__6_,
         mem_stage_inst_dmem_ram_80__7_, mem_stage_inst_dmem_ram_80__8_,
         mem_stage_inst_dmem_ram_80__9_, mem_stage_inst_dmem_ram_80__10_,
         mem_stage_inst_dmem_ram_80__11_, mem_stage_inst_dmem_ram_80__12_,
         mem_stage_inst_dmem_ram_80__13_, mem_stage_inst_dmem_ram_80__14_,
         mem_stage_inst_dmem_ram_80__15_, mem_stage_inst_dmem_ram_81__0_,
         mem_stage_inst_dmem_ram_81__1_, mem_stage_inst_dmem_ram_81__2_,
         mem_stage_inst_dmem_ram_81__3_, mem_stage_inst_dmem_ram_81__4_,
         mem_stage_inst_dmem_ram_81__5_, mem_stage_inst_dmem_ram_81__6_,
         mem_stage_inst_dmem_ram_81__7_, mem_stage_inst_dmem_ram_81__8_,
         mem_stage_inst_dmem_ram_81__9_, mem_stage_inst_dmem_ram_81__10_,
         mem_stage_inst_dmem_ram_81__11_, mem_stage_inst_dmem_ram_81__12_,
         mem_stage_inst_dmem_ram_81__13_, mem_stage_inst_dmem_ram_81__14_,
         mem_stage_inst_dmem_ram_81__15_, mem_stage_inst_dmem_ram_82__0_,
         mem_stage_inst_dmem_ram_82__1_, mem_stage_inst_dmem_ram_82__2_,
         mem_stage_inst_dmem_ram_82__3_, mem_stage_inst_dmem_ram_82__4_,
         mem_stage_inst_dmem_ram_82__5_, mem_stage_inst_dmem_ram_82__6_,
         mem_stage_inst_dmem_ram_82__7_, mem_stage_inst_dmem_ram_82__8_,
         mem_stage_inst_dmem_ram_82__9_, mem_stage_inst_dmem_ram_82__10_,
         mem_stage_inst_dmem_ram_82__11_, mem_stage_inst_dmem_ram_82__12_,
         mem_stage_inst_dmem_ram_82__13_, mem_stage_inst_dmem_ram_82__14_,
         mem_stage_inst_dmem_ram_82__15_, mem_stage_inst_dmem_ram_83__0_,
         mem_stage_inst_dmem_ram_83__1_, mem_stage_inst_dmem_ram_83__2_,
         mem_stage_inst_dmem_ram_83__3_, mem_stage_inst_dmem_ram_83__4_,
         mem_stage_inst_dmem_ram_83__5_, mem_stage_inst_dmem_ram_83__6_,
         mem_stage_inst_dmem_ram_83__7_, mem_stage_inst_dmem_ram_83__8_,
         mem_stage_inst_dmem_ram_83__9_, mem_stage_inst_dmem_ram_83__10_,
         mem_stage_inst_dmem_ram_83__11_, mem_stage_inst_dmem_ram_83__12_,
         mem_stage_inst_dmem_ram_83__13_, mem_stage_inst_dmem_ram_83__14_,
         mem_stage_inst_dmem_ram_83__15_, mem_stage_inst_dmem_ram_84__0_,
         mem_stage_inst_dmem_ram_84__1_, mem_stage_inst_dmem_ram_84__2_,
         mem_stage_inst_dmem_ram_84__3_, mem_stage_inst_dmem_ram_84__4_,
         mem_stage_inst_dmem_ram_84__5_, mem_stage_inst_dmem_ram_84__6_,
         mem_stage_inst_dmem_ram_84__7_, mem_stage_inst_dmem_ram_84__8_,
         mem_stage_inst_dmem_ram_84__9_, mem_stage_inst_dmem_ram_84__10_,
         mem_stage_inst_dmem_ram_84__11_, mem_stage_inst_dmem_ram_84__12_,
         mem_stage_inst_dmem_ram_84__13_, mem_stage_inst_dmem_ram_84__14_,
         mem_stage_inst_dmem_ram_84__15_, mem_stage_inst_dmem_ram_85__0_,
         mem_stage_inst_dmem_ram_85__1_, mem_stage_inst_dmem_ram_85__2_,
         mem_stage_inst_dmem_ram_85__3_, mem_stage_inst_dmem_ram_85__4_,
         mem_stage_inst_dmem_ram_85__5_, mem_stage_inst_dmem_ram_85__6_,
         mem_stage_inst_dmem_ram_85__7_, mem_stage_inst_dmem_ram_85__8_,
         mem_stage_inst_dmem_ram_85__9_, mem_stage_inst_dmem_ram_85__10_,
         mem_stage_inst_dmem_ram_85__11_, mem_stage_inst_dmem_ram_85__12_,
         mem_stage_inst_dmem_ram_85__13_, mem_stage_inst_dmem_ram_85__14_,
         mem_stage_inst_dmem_ram_85__15_, mem_stage_inst_dmem_ram_86__0_,
         mem_stage_inst_dmem_ram_86__1_, mem_stage_inst_dmem_ram_86__2_,
         mem_stage_inst_dmem_ram_86__3_, mem_stage_inst_dmem_ram_86__4_,
         mem_stage_inst_dmem_ram_86__5_, mem_stage_inst_dmem_ram_86__6_,
         mem_stage_inst_dmem_ram_86__7_, mem_stage_inst_dmem_ram_86__8_,
         mem_stage_inst_dmem_ram_86__9_, mem_stage_inst_dmem_ram_86__10_,
         mem_stage_inst_dmem_ram_86__11_, mem_stage_inst_dmem_ram_86__12_,
         mem_stage_inst_dmem_ram_86__13_, mem_stage_inst_dmem_ram_86__14_,
         mem_stage_inst_dmem_ram_86__15_, mem_stage_inst_dmem_ram_87__0_,
         mem_stage_inst_dmem_ram_87__1_, mem_stage_inst_dmem_ram_87__2_,
         mem_stage_inst_dmem_ram_87__3_, mem_stage_inst_dmem_ram_87__4_,
         mem_stage_inst_dmem_ram_87__5_, mem_stage_inst_dmem_ram_87__6_,
         mem_stage_inst_dmem_ram_87__7_, mem_stage_inst_dmem_ram_87__8_,
         mem_stage_inst_dmem_ram_87__9_, mem_stage_inst_dmem_ram_87__10_,
         mem_stage_inst_dmem_ram_87__11_, mem_stage_inst_dmem_ram_87__12_,
         mem_stage_inst_dmem_ram_87__13_, mem_stage_inst_dmem_ram_87__14_,
         mem_stage_inst_dmem_ram_87__15_, mem_stage_inst_dmem_ram_88__0_,
         mem_stage_inst_dmem_ram_88__1_, mem_stage_inst_dmem_ram_88__2_,
         mem_stage_inst_dmem_ram_88__3_, mem_stage_inst_dmem_ram_88__4_,
         mem_stage_inst_dmem_ram_88__5_, mem_stage_inst_dmem_ram_88__6_,
         mem_stage_inst_dmem_ram_88__7_, mem_stage_inst_dmem_ram_88__8_,
         mem_stage_inst_dmem_ram_88__9_, mem_stage_inst_dmem_ram_88__10_,
         mem_stage_inst_dmem_ram_88__11_, mem_stage_inst_dmem_ram_88__12_,
         mem_stage_inst_dmem_ram_88__13_, mem_stage_inst_dmem_ram_88__14_,
         mem_stage_inst_dmem_ram_88__15_, mem_stage_inst_dmem_ram_89__0_,
         mem_stage_inst_dmem_ram_89__1_, mem_stage_inst_dmem_ram_89__2_,
         mem_stage_inst_dmem_ram_89__3_, mem_stage_inst_dmem_ram_89__4_,
         mem_stage_inst_dmem_ram_89__5_, mem_stage_inst_dmem_ram_89__6_,
         mem_stage_inst_dmem_ram_89__7_, mem_stage_inst_dmem_ram_89__8_,
         mem_stage_inst_dmem_ram_89__9_, mem_stage_inst_dmem_ram_89__10_,
         mem_stage_inst_dmem_ram_89__11_, mem_stage_inst_dmem_ram_89__12_,
         mem_stage_inst_dmem_ram_89__13_, mem_stage_inst_dmem_ram_89__14_,
         mem_stage_inst_dmem_ram_89__15_, mem_stage_inst_dmem_ram_90__0_,
         mem_stage_inst_dmem_ram_90__1_, mem_stage_inst_dmem_ram_90__2_,
         mem_stage_inst_dmem_ram_90__3_, mem_stage_inst_dmem_ram_90__4_,
         mem_stage_inst_dmem_ram_90__5_, mem_stage_inst_dmem_ram_90__6_,
         mem_stage_inst_dmem_ram_90__7_, mem_stage_inst_dmem_ram_90__8_,
         mem_stage_inst_dmem_ram_90__9_, mem_stage_inst_dmem_ram_90__10_,
         mem_stage_inst_dmem_ram_90__11_, mem_stage_inst_dmem_ram_90__12_,
         mem_stage_inst_dmem_ram_90__13_, mem_stage_inst_dmem_ram_90__14_,
         mem_stage_inst_dmem_ram_90__15_, mem_stage_inst_dmem_ram_91__0_,
         mem_stage_inst_dmem_ram_91__1_, mem_stage_inst_dmem_ram_91__2_,
         mem_stage_inst_dmem_ram_91__3_, mem_stage_inst_dmem_ram_91__4_,
         mem_stage_inst_dmem_ram_91__5_, mem_stage_inst_dmem_ram_91__6_,
         mem_stage_inst_dmem_ram_91__7_, mem_stage_inst_dmem_ram_91__8_,
         mem_stage_inst_dmem_ram_91__9_, mem_stage_inst_dmem_ram_91__10_,
         mem_stage_inst_dmem_ram_91__11_, mem_stage_inst_dmem_ram_91__12_,
         mem_stage_inst_dmem_ram_91__13_, mem_stage_inst_dmem_ram_91__14_,
         mem_stage_inst_dmem_ram_91__15_, mem_stage_inst_dmem_ram_92__0_,
         mem_stage_inst_dmem_ram_92__1_, mem_stage_inst_dmem_ram_92__2_,
         mem_stage_inst_dmem_ram_92__3_, mem_stage_inst_dmem_ram_92__4_,
         mem_stage_inst_dmem_ram_92__5_, mem_stage_inst_dmem_ram_92__6_,
         mem_stage_inst_dmem_ram_92__7_, mem_stage_inst_dmem_ram_92__8_,
         mem_stage_inst_dmem_ram_92__9_, mem_stage_inst_dmem_ram_92__10_,
         mem_stage_inst_dmem_ram_92__11_, mem_stage_inst_dmem_ram_92__12_,
         mem_stage_inst_dmem_ram_92__13_, mem_stage_inst_dmem_ram_92__14_,
         mem_stage_inst_dmem_ram_92__15_, mem_stage_inst_dmem_ram_93__0_,
         mem_stage_inst_dmem_ram_93__1_, mem_stage_inst_dmem_ram_93__2_,
         mem_stage_inst_dmem_ram_93__3_, mem_stage_inst_dmem_ram_93__4_,
         mem_stage_inst_dmem_ram_93__5_, mem_stage_inst_dmem_ram_93__6_,
         mem_stage_inst_dmem_ram_93__7_, mem_stage_inst_dmem_ram_93__8_,
         mem_stage_inst_dmem_ram_93__9_, mem_stage_inst_dmem_ram_93__10_,
         mem_stage_inst_dmem_ram_93__11_, mem_stage_inst_dmem_ram_93__12_,
         mem_stage_inst_dmem_ram_93__13_, mem_stage_inst_dmem_ram_93__14_,
         mem_stage_inst_dmem_ram_93__15_, mem_stage_inst_dmem_ram_94__0_,
         mem_stage_inst_dmem_ram_94__1_, mem_stage_inst_dmem_ram_94__2_,
         mem_stage_inst_dmem_ram_94__3_, mem_stage_inst_dmem_ram_94__4_,
         mem_stage_inst_dmem_ram_94__5_, mem_stage_inst_dmem_ram_94__6_,
         mem_stage_inst_dmem_ram_94__7_, mem_stage_inst_dmem_ram_94__8_,
         mem_stage_inst_dmem_ram_94__9_, mem_stage_inst_dmem_ram_94__10_,
         mem_stage_inst_dmem_ram_94__11_, mem_stage_inst_dmem_ram_94__12_,
         mem_stage_inst_dmem_ram_94__13_, mem_stage_inst_dmem_ram_94__14_,
         mem_stage_inst_dmem_ram_94__15_, mem_stage_inst_dmem_ram_95__0_,
         mem_stage_inst_dmem_ram_95__1_, mem_stage_inst_dmem_ram_95__2_,
         mem_stage_inst_dmem_ram_95__3_, mem_stage_inst_dmem_ram_95__4_,
         mem_stage_inst_dmem_ram_95__5_, mem_stage_inst_dmem_ram_95__6_,
         mem_stage_inst_dmem_ram_95__7_, mem_stage_inst_dmem_ram_95__8_,
         mem_stage_inst_dmem_ram_95__9_, mem_stage_inst_dmem_ram_95__10_,
         mem_stage_inst_dmem_ram_95__11_, mem_stage_inst_dmem_ram_95__12_,
         mem_stage_inst_dmem_ram_95__13_, mem_stage_inst_dmem_ram_95__14_,
         mem_stage_inst_dmem_ram_95__15_, mem_stage_inst_dmem_ram_32__0_,
         mem_stage_inst_dmem_ram_32__1_, mem_stage_inst_dmem_ram_32__2_,
         mem_stage_inst_dmem_ram_32__3_, mem_stage_inst_dmem_ram_32__4_,
         mem_stage_inst_dmem_ram_32__5_, mem_stage_inst_dmem_ram_32__6_,
         mem_stage_inst_dmem_ram_32__7_, mem_stage_inst_dmem_ram_32__8_,
         mem_stage_inst_dmem_ram_32__9_, mem_stage_inst_dmem_ram_32__10_,
         mem_stage_inst_dmem_ram_32__11_, mem_stage_inst_dmem_ram_32__12_,
         mem_stage_inst_dmem_ram_32__13_, mem_stage_inst_dmem_ram_32__14_,
         mem_stage_inst_dmem_ram_32__15_, mem_stage_inst_dmem_ram_33__0_,
         mem_stage_inst_dmem_ram_33__1_, mem_stage_inst_dmem_ram_33__2_,
         mem_stage_inst_dmem_ram_33__3_, mem_stage_inst_dmem_ram_33__4_,
         mem_stage_inst_dmem_ram_33__5_, mem_stage_inst_dmem_ram_33__6_,
         mem_stage_inst_dmem_ram_33__7_, mem_stage_inst_dmem_ram_33__8_,
         mem_stage_inst_dmem_ram_33__9_, mem_stage_inst_dmem_ram_33__10_,
         mem_stage_inst_dmem_ram_33__11_, mem_stage_inst_dmem_ram_33__12_,
         mem_stage_inst_dmem_ram_33__13_, mem_stage_inst_dmem_ram_33__14_,
         mem_stage_inst_dmem_ram_33__15_, mem_stage_inst_dmem_ram_34__0_,
         mem_stage_inst_dmem_ram_34__1_, mem_stage_inst_dmem_ram_34__2_,
         mem_stage_inst_dmem_ram_34__3_, mem_stage_inst_dmem_ram_34__4_,
         mem_stage_inst_dmem_ram_34__5_, mem_stage_inst_dmem_ram_34__6_,
         mem_stage_inst_dmem_ram_34__7_, mem_stage_inst_dmem_ram_34__8_,
         mem_stage_inst_dmem_ram_34__9_, mem_stage_inst_dmem_ram_34__10_,
         mem_stage_inst_dmem_ram_34__11_, mem_stage_inst_dmem_ram_34__12_,
         mem_stage_inst_dmem_ram_34__13_, mem_stage_inst_dmem_ram_34__14_,
         mem_stage_inst_dmem_ram_34__15_, mem_stage_inst_dmem_ram_35__0_,
         mem_stage_inst_dmem_ram_35__1_, mem_stage_inst_dmem_ram_35__2_,
         mem_stage_inst_dmem_ram_35__3_, mem_stage_inst_dmem_ram_35__4_,
         mem_stage_inst_dmem_ram_35__5_, mem_stage_inst_dmem_ram_35__6_,
         mem_stage_inst_dmem_ram_35__7_, mem_stage_inst_dmem_ram_35__8_,
         mem_stage_inst_dmem_ram_35__9_, mem_stage_inst_dmem_ram_35__10_,
         mem_stage_inst_dmem_ram_35__11_, mem_stage_inst_dmem_ram_35__12_,
         mem_stage_inst_dmem_ram_35__13_, mem_stage_inst_dmem_ram_35__14_,
         mem_stage_inst_dmem_ram_35__15_, mem_stage_inst_dmem_ram_36__0_,
         mem_stage_inst_dmem_ram_36__1_, mem_stage_inst_dmem_ram_36__2_,
         mem_stage_inst_dmem_ram_36__3_, mem_stage_inst_dmem_ram_36__4_,
         mem_stage_inst_dmem_ram_36__5_, mem_stage_inst_dmem_ram_36__6_,
         mem_stage_inst_dmem_ram_36__7_, mem_stage_inst_dmem_ram_36__8_,
         mem_stage_inst_dmem_ram_36__9_, mem_stage_inst_dmem_ram_36__10_,
         mem_stage_inst_dmem_ram_36__11_, mem_stage_inst_dmem_ram_36__12_,
         mem_stage_inst_dmem_ram_36__13_, mem_stage_inst_dmem_ram_36__14_,
         mem_stage_inst_dmem_ram_36__15_, mem_stage_inst_dmem_ram_37__0_,
         mem_stage_inst_dmem_ram_37__1_, mem_stage_inst_dmem_ram_37__2_,
         mem_stage_inst_dmem_ram_37__3_, mem_stage_inst_dmem_ram_37__4_,
         mem_stage_inst_dmem_ram_37__5_, mem_stage_inst_dmem_ram_37__6_,
         mem_stage_inst_dmem_ram_37__7_, mem_stage_inst_dmem_ram_37__8_,
         mem_stage_inst_dmem_ram_37__9_, mem_stage_inst_dmem_ram_37__10_,
         mem_stage_inst_dmem_ram_37__11_, mem_stage_inst_dmem_ram_37__12_,
         mem_stage_inst_dmem_ram_37__13_, mem_stage_inst_dmem_ram_37__14_,
         mem_stage_inst_dmem_ram_37__15_, mem_stage_inst_dmem_ram_38__0_,
         mem_stage_inst_dmem_ram_38__1_, mem_stage_inst_dmem_ram_38__2_,
         mem_stage_inst_dmem_ram_38__3_, mem_stage_inst_dmem_ram_38__4_,
         mem_stage_inst_dmem_ram_38__5_, mem_stage_inst_dmem_ram_38__6_,
         mem_stage_inst_dmem_ram_38__7_, mem_stage_inst_dmem_ram_38__8_,
         mem_stage_inst_dmem_ram_38__9_, mem_stage_inst_dmem_ram_38__10_,
         mem_stage_inst_dmem_ram_38__11_, mem_stage_inst_dmem_ram_38__12_,
         mem_stage_inst_dmem_ram_38__13_, mem_stage_inst_dmem_ram_38__14_,
         mem_stage_inst_dmem_ram_38__15_, mem_stage_inst_dmem_ram_39__0_,
         mem_stage_inst_dmem_ram_39__1_, mem_stage_inst_dmem_ram_39__2_,
         mem_stage_inst_dmem_ram_39__3_, mem_stage_inst_dmem_ram_39__4_,
         mem_stage_inst_dmem_ram_39__5_, mem_stage_inst_dmem_ram_39__6_,
         mem_stage_inst_dmem_ram_39__7_, mem_stage_inst_dmem_ram_39__8_,
         mem_stage_inst_dmem_ram_39__9_, mem_stage_inst_dmem_ram_39__10_,
         mem_stage_inst_dmem_ram_39__11_, mem_stage_inst_dmem_ram_39__12_,
         mem_stage_inst_dmem_ram_39__13_, mem_stage_inst_dmem_ram_39__14_,
         mem_stage_inst_dmem_ram_39__15_, mem_stage_inst_dmem_ram_40__0_,
         mem_stage_inst_dmem_ram_40__1_, mem_stage_inst_dmem_ram_40__2_,
         mem_stage_inst_dmem_ram_40__3_, mem_stage_inst_dmem_ram_40__4_,
         mem_stage_inst_dmem_ram_40__5_, mem_stage_inst_dmem_ram_40__6_,
         mem_stage_inst_dmem_ram_40__7_, mem_stage_inst_dmem_ram_40__8_,
         mem_stage_inst_dmem_ram_40__9_, mem_stage_inst_dmem_ram_40__10_,
         mem_stage_inst_dmem_ram_40__11_, mem_stage_inst_dmem_ram_40__12_,
         mem_stage_inst_dmem_ram_40__13_, mem_stage_inst_dmem_ram_40__14_,
         mem_stage_inst_dmem_ram_40__15_, mem_stage_inst_dmem_ram_41__0_,
         mem_stage_inst_dmem_ram_41__1_, mem_stage_inst_dmem_ram_41__2_,
         mem_stage_inst_dmem_ram_41__3_, mem_stage_inst_dmem_ram_41__4_,
         mem_stage_inst_dmem_ram_41__5_, mem_stage_inst_dmem_ram_41__6_,
         mem_stage_inst_dmem_ram_41__7_, mem_stage_inst_dmem_ram_41__8_,
         mem_stage_inst_dmem_ram_41__9_, mem_stage_inst_dmem_ram_41__10_,
         mem_stage_inst_dmem_ram_41__11_, mem_stage_inst_dmem_ram_41__12_,
         mem_stage_inst_dmem_ram_41__13_, mem_stage_inst_dmem_ram_41__14_,
         mem_stage_inst_dmem_ram_41__15_, mem_stage_inst_dmem_ram_42__0_,
         mem_stage_inst_dmem_ram_42__1_, mem_stage_inst_dmem_ram_42__2_,
         mem_stage_inst_dmem_ram_42__3_, mem_stage_inst_dmem_ram_42__4_,
         mem_stage_inst_dmem_ram_42__5_, mem_stage_inst_dmem_ram_42__6_,
         mem_stage_inst_dmem_ram_42__7_, mem_stage_inst_dmem_ram_42__8_,
         mem_stage_inst_dmem_ram_42__9_, mem_stage_inst_dmem_ram_42__10_,
         mem_stage_inst_dmem_ram_42__11_, mem_stage_inst_dmem_ram_42__12_,
         mem_stage_inst_dmem_ram_42__13_, mem_stage_inst_dmem_ram_42__14_,
         mem_stage_inst_dmem_ram_42__15_, mem_stage_inst_dmem_ram_43__0_,
         mem_stage_inst_dmem_ram_43__1_, mem_stage_inst_dmem_ram_43__2_,
         mem_stage_inst_dmem_ram_43__3_, mem_stage_inst_dmem_ram_43__4_,
         mem_stage_inst_dmem_ram_43__5_, mem_stage_inst_dmem_ram_43__6_,
         mem_stage_inst_dmem_ram_43__7_, mem_stage_inst_dmem_ram_43__8_,
         mem_stage_inst_dmem_ram_43__9_, mem_stage_inst_dmem_ram_43__10_,
         mem_stage_inst_dmem_ram_43__11_, mem_stage_inst_dmem_ram_43__12_,
         mem_stage_inst_dmem_ram_43__13_, mem_stage_inst_dmem_ram_43__14_,
         mem_stage_inst_dmem_ram_43__15_, mem_stage_inst_dmem_ram_44__0_,
         mem_stage_inst_dmem_ram_44__1_, mem_stage_inst_dmem_ram_44__2_,
         mem_stage_inst_dmem_ram_44__3_, mem_stage_inst_dmem_ram_44__4_,
         mem_stage_inst_dmem_ram_44__5_, mem_stage_inst_dmem_ram_44__6_,
         mem_stage_inst_dmem_ram_44__7_, mem_stage_inst_dmem_ram_44__8_,
         mem_stage_inst_dmem_ram_44__9_, mem_stage_inst_dmem_ram_44__10_,
         mem_stage_inst_dmem_ram_44__11_, mem_stage_inst_dmem_ram_44__12_,
         mem_stage_inst_dmem_ram_44__13_, mem_stage_inst_dmem_ram_44__14_,
         mem_stage_inst_dmem_ram_44__15_, mem_stage_inst_dmem_ram_45__0_,
         mem_stage_inst_dmem_ram_45__1_, mem_stage_inst_dmem_ram_45__2_,
         mem_stage_inst_dmem_ram_45__3_, mem_stage_inst_dmem_ram_45__4_,
         mem_stage_inst_dmem_ram_45__5_, mem_stage_inst_dmem_ram_45__6_,
         mem_stage_inst_dmem_ram_45__7_, mem_stage_inst_dmem_ram_45__8_,
         mem_stage_inst_dmem_ram_45__9_, mem_stage_inst_dmem_ram_45__10_,
         mem_stage_inst_dmem_ram_45__11_, mem_stage_inst_dmem_ram_45__12_,
         mem_stage_inst_dmem_ram_45__13_, mem_stage_inst_dmem_ram_45__14_,
         mem_stage_inst_dmem_ram_45__15_, mem_stage_inst_dmem_ram_46__0_,
         mem_stage_inst_dmem_ram_46__1_, mem_stage_inst_dmem_ram_46__2_,
         mem_stage_inst_dmem_ram_46__3_, mem_stage_inst_dmem_ram_46__4_,
         mem_stage_inst_dmem_ram_46__5_, mem_stage_inst_dmem_ram_46__6_,
         mem_stage_inst_dmem_ram_46__7_, mem_stage_inst_dmem_ram_46__8_,
         mem_stage_inst_dmem_ram_46__9_, mem_stage_inst_dmem_ram_46__10_,
         mem_stage_inst_dmem_ram_46__11_, mem_stage_inst_dmem_ram_46__12_,
         mem_stage_inst_dmem_ram_46__13_, mem_stage_inst_dmem_ram_46__14_,
         mem_stage_inst_dmem_ram_46__15_, mem_stage_inst_dmem_ram_47__0_,
         mem_stage_inst_dmem_ram_47__1_, mem_stage_inst_dmem_ram_47__2_,
         mem_stage_inst_dmem_ram_47__3_, mem_stage_inst_dmem_ram_47__4_,
         mem_stage_inst_dmem_ram_47__5_, mem_stage_inst_dmem_ram_47__6_,
         mem_stage_inst_dmem_ram_47__7_, mem_stage_inst_dmem_ram_47__8_,
         mem_stage_inst_dmem_ram_47__9_, mem_stage_inst_dmem_ram_47__10_,
         mem_stage_inst_dmem_ram_47__11_, mem_stage_inst_dmem_ram_47__12_,
         mem_stage_inst_dmem_ram_47__13_, mem_stage_inst_dmem_ram_47__14_,
         mem_stage_inst_dmem_ram_47__15_, mem_stage_inst_dmem_ram_48__0_,
         mem_stage_inst_dmem_ram_48__1_, mem_stage_inst_dmem_ram_48__2_,
         mem_stage_inst_dmem_ram_48__3_, mem_stage_inst_dmem_ram_48__4_,
         mem_stage_inst_dmem_ram_48__5_, mem_stage_inst_dmem_ram_48__6_,
         mem_stage_inst_dmem_ram_48__7_, mem_stage_inst_dmem_ram_48__8_,
         mem_stage_inst_dmem_ram_48__9_, mem_stage_inst_dmem_ram_48__10_,
         mem_stage_inst_dmem_ram_48__11_, mem_stage_inst_dmem_ram_48__12_,
         mem_stage_inst_dmem_ram_48__13_, mem_stage_inst_dmem_ram_48__14_,
         mem_stage_inst_dmem_ram_48__15_, mem_stage_inst_dmem_ram_49__0_,
         mem_stage_inst_dmem_ram_49__1_, mem_stage_inst_dmem_ram_49__2_,
         mem_stage_inst_dmem_ram_49__3_, mem_stage_inst_dmem_ram_49__4_,
         mem_stage_inst_dmem_ram_49__5_, mem_stage_inst_dmem_ram_49__6_,
         mem_stage_inst_dmem_ram_49__7_, mem_stage_inst_dmem_ram_49__8_,
         mem_stage_inst_dmem_ram_49__9_, mem_stage_inst_dmem_ram_49__10_,
         mem_stage_inst_dmem_ram_49__11_, mem_stage_inst_dmem_ram_49__12_,
         mem_stage_inst_dmem_ram_49__13_, mem_stage_inst_dmem_ram_49__14_,
         mem_stage_inst_dmem_ram_49__15_, mem_stage_inst_dmem_ram_50__0_,
         mem_stage_inst_dmem_ram_50__1_, mem_stage_inst_dmem_ram_50__2_,
         mem_stage_inst_dmem_ram_50__3_, mem_stage_inst_dmem_ram_50__4_,
         mem_stage_inst_dmem_ram_50__5_, mem_stage_inst_dmem_ram_50__6_,
         mem_stage_inst_dmem_ram_50__7_, mem_stage_inst_dmem_ram_50__8_,
         mem_stage_inst_dmem_ram_50__9_, mem_stage_inst_dmem_ram_50__10_,
         mem_stage_inst_dmem_ram_50__11_, mem_stage_inst_dmem_ram_50__12_,
         mem_stage_inst_dmem_ram_50__13_, mem_stage_inst_dmem_ram_50__14_,
         mem_stage_inst_dmem_ram_50__15_, mem_stage_inst_dmem_ram_51__0_,
         mem_stage_inst_dmem_ram_51__1_, mem_stage_inst_dmem_ram_51__2_,
         mem_stage_inst_dmem_ram_51__3_, mem_stage_inst_dmem_ram_51__4_,
         mem_stage_inst_dmem_ram_51__5_, mem_stage_inst_dmem_ram_51__6_,
         mem_stage_inst_dmem_ram_51__7_, mem_stage_inst_dmem_ram_51__8_,
         mem_stage_inst_dmem_ram_51__9_, mem_stage_inst_dmem_ram_51__10_,
         mem_stage_inst_dmem_ram_51__11_, mem_stage_inst_dmem_ram_51__12_,
         mem_stage_inst_dmem_ram_51__13_, mem_stage_inst_dmem_ram_51__14_,
         mem_stage_inst_dmem_ram_51__15_, mem_stage_inst_dmem_ram_52__0_,
         mem_stage_inst_dmem_ram_52__1_, mem_stage_inst_dmem_ram_52__2_,
         mem_stage_inst_dmem_ram_52__3_, mem_stage_inst_dmem_ram_52__4_,
         mem_stage_inst_dmem_ram_52__5_, mem_stage_inst_dmem_ram_52__6_,
         mem_stage_inst_dmem_ram_52__7_, mem_stage_inst_dmem_ram_52__8_,
         mem_stage_inst_dmem_ram_52__9_, mem_stage_inst_dmem_ram_52__10_,
         mem_stage_inst_dmem_ram_52__11_, mem_stage_inst_dmem_ram_52__12_,
         mem_stage_inst_dmem_ram_52__13_, mem_stage_inst_dmem_ram_52__14_,
         mem_stage_inst_dmem_ram_52__15_, mem_stage_inst_dmem_ram_53__0_,
         mem_stage_inst_dmem_ram_53__1_, mem_stage_inst_dmem_ram_53__2_,
         mem_stage_inst_dmem_ram_53__3_, mem_stage_inst_dmem_ram_53__4_,
         mem_stage_inst_dmem_ram_53__5_, mem_stage_inst_dmem_ram_53__6_,
         mem_stage_inst_dmem_ram_53__7_, mem_stage_inst_dmem_ram_53__8_,
         mem_stage_inst_dmem_ram_53__9_, mem_stage_inst_dmem_ram_53__10_,
         mem_stage_inst_dmem_ram_53__11_, mem_stage_inst_dmem_ram_53__12_,
         mem_stage_inst_dmem_ram_53__13_, mem_stage_inst_dmem_ram_53__14_,
         mem_stage_inst_dmem_ram_53__15_, mem_stage_inst_dmem_ram_54__0_,
         mem_stage_inst_dmem_ram_54__1_, mem_stage_inst_dmem_ram_54__2_,
         mem_stage_inst_dmem_ram_54__3_, mem_stage_inst_dmem_ram_54__4_,
         mem_stage_inst_dmem_ram_54__5_, mem_stage_inst_dmem_ram_54__6_,
         mem_stage_inst_dmem_ram_54__7_, mem_stage_inst_dmem_ram_54__8_,
         mem_stage_inst_dmem_ram_54__9_, mem_stage_inst_dmem_ram_54__10_,
         mem_stage_inst_dmem_ram_54__11_, mem_stage_inst_dmem_ram_54__12_,
         mem_stage_inst_dmem_ram_54__13_, mem_stage_inst_dmem_ram_54__14_,
         mem_stage_inst_dmem_ram_54__15_, mem_stage_inst_dmem_ram_55__0_,
         mem_stage_inst_dmem_ram_55__1_, mem_stage_inst_dmem_ram_55__2_,
         mem_stage_inst_dmem_ram_55__3_, mem_stage_inst_dmem_ram_55__4_,
         mem_stage_inst_dmem_ram_55__5_, mem_stage_inst_dmem_ram_55__6_,
         mem_stage_inst_dmem_ram_55__7_, mem_stage_inst_dmem_ram_55__8_,
         mem_stage_inst_dmem_ram_55__9_, mem_stage_inst_dmem_ram_55__10_,
         mem_stage_inst_dmem_ram_55__11_, mem_stage_inst_dmem_ram_55__12_,
         mem_stage_inst_dmem_ram_55__13_, mem_stage_inst_dmem_ram_55__14_,
         mem_stage_inst_dmem_ram_55__15_, mem_stage_inst_dmem_ram_56__0_,
         mem_stage_inst_dmem_ram_56__1_, mem_stage_inst_dmem_ram_56__2_,
         mem_stage_inst_dmem_ram_56__3_, mem_stage_inst_dmem_ram_56__4_,
         mem_stage_inst_dmem_ram_56__5_, mem_stage_inst_dmem_ram_56__6_,
         mem_stage_inst_dmem_ram_56__7_, mem_stage_inst_dmem_ram_56__8_,
         mem_stage_inst_dmem_ram_56__9_, mem_stage_inst_dmem_ram_56__10_,
         mem_stage_inst_dmem_ram_56__11_, mem_stage_inst_dmem_ram_56__12_,
         mem_stage_inst_dmem_ram_56__13_, mem_stage_inst_dmem_ram_56__14_,
         mem_stage_inst_dmem_ram_56__15_, mem_stage_inst_dmem_ram_57__0_,
         mem_stage_inst_dmem_ram_57__1_, mem_stage_inst_dmem_ram_57__2_,
         mem_stage_inst_dmem_ram_57__3_, mem_stage_inst_dmem_ram_57__4_,
         mem_stage_inst_dmem_ram_57__5_, mem_stage_inst_dmem_ram_57__6_,
         mem_stage_inst_dmem_ram_57__7_, mem_stage_inst_dmem_ram_57__8_,
         mem_stage_inst_dmem_ram_57__9_, mem_stage_inst_dmem_ram_57__10_,
         mem_stage_inst_dmem_ram_57__11_, mem_stage_inst_dmem_ram_57__12_,
         mem_stage_inst_dmem_ram_57__13_, mem_stage_inst_dmem_ram_57__14_,
         mem_stage_inst_dmem_ram_57__15_, mem_stage_inst_dmem_ram_58__0_,
         mem_stage_inst_dmem_ram_58__1_, mem_stage_inst_dmem_ram_58__2_,
         mem_stage_inst_dmem_ram_58__3_, mem_stage_inst_dmem_ram_58__4_,
         mem_stage_inst_dmem_ram_58__5_, mem_stage_inst_dmem_ram_58__6_,
         mem_stage_inst_dmem_ram_58__7_, mem_stage_inst_dmem_ram_58__8_,
         mem_stage_inst_dmem_ram_58__9_, mem_stage_inst_dmem_ram_58__10_,
         mem_stage_inst_dmem_ram_58__11_, mem_stage_inst_dmem_ram_58__12_,
         mem_stage_inst_dmem_ram_58__13_, mem_stage_inst_dmem_ram_58__14_,
         mem_stage_inst_dmem_ram_58__15_, mem_stage_inst_dmem_ram_59__0_,
         mem_stage_inst_dmem_ram_59__1_, mem_stage_inst_dmem_ram_59__2_,
         mem_stage_inst_dmem_ram_59__3_, mem_stage_inst_dmem_ram_59__4_,
         mem_stage_inst_dmem_ram_59__5_, mem_stage_inst_dmem_ram_59__6_,
         mem_stage_inst_dmem_ram_59__7_, mem_stage_inst_dmem_ram_59__8_,
         mem_stage_inst_dmem_ram_59__9_, mem_stage_inst_dmem_ram_59__10_,
         mem_stage_inst_dmem_ram_59__11_, mem_stage_inst_dmem_ram_59__12_,
         mem_stage_inst_dmem_ram_59__13_, mem_stage_inst_dmem_ram_59__14_,
         mem_stage_inst_dmem_ram_59__15_, mem_stage_inst_dmem_ram_60__0_,
         mem_stage_inst_dmem_ram_60__1_, mem_stage_inst_dmem_ram_60__2_,
         mem_stage_inst_dmem_ram_60__3_, mem_stage_inst_dmem_ram_60__4_,
         mem_stage_inst_dmem_ram_60__5_, mem_stage_inst_dmem_ram_60__6_,
         mem_stage_inst_dmem_ram_60__7_, mem_stage_inst_dmem_ram_60__8_,
         mem_stage_inst_dmem_ram_60__9_, mem_stage_inst_dmem_ram_60__10_,
         mem_stage_inst_dmem_ram_60__11_, mem_stage_inst_dmem_ram_60__12_,
         mem_stage_inst_dmem_ram_60__13_, mem_stage_inst_dmem_ram_60__14_,
         mem_stage_inst_dmem_ram_60__15_, mem_stage_inst_dmem_ram_61__0_,
         mem_stage_inst_dmem_ram_61__1_, mem_stage_inst_dmem_ram_61__2_,
         mem_stage_inst_dmem_ram_61__3_, mem_stage_inst_dmem_ram_61__4_,
         mem_stage_inst_dmem_ram_61__5_, mem_stage_inst_dmem_ram_61__6_,
         mem_stage_inst_dmem_ram_61__7_, mem_stage_inst_dmem_ram_61__8_,
         mem_stage_inst_dmem_ram_61__9_, mem_stage_inst_dmem_ram_61__10_,
         mem_stage_inst_dmem_ram_61__11_, mem_stage_inst_dmem_ram_61__12_,
         mem_stage_inst_dmem_ram_61__13_, mem_stage_inst_dmem_ram_61__14_,
         mem_stage_inst_dmem_ram_61__15_, mem_stage_inst_dmem_ram_62__0_,
         mem_stage_inst_dmem_ram_62__1_, mem_stage_inst_dmem_ram_62__2_,
         mem_stage_inst_dmem_ram_62__3_, mem_stage_inst_dmem_ram_62__4_,
         mem_stage_inst_dmem_ram_62__5_, mem_stage_inst_dmem_ram_62__6_,
         mem_stage_inst_dmem_ram_62__7_, mem_stage_inst_dmem_ram_62__8_,
         mem_stage_inst_dmem_ram_62__9_, mem_stage_inst_dmem_ram_62__10_,
         mem_stage_inst_dmem_ram_62__11_, mem_stage_inst_dmem_ram_62__12_,
         mem_stage_inst_dmem_ram_62__13_, mem_stage_inst_dmem_ram_62__14_,
         mem_stage_inst_dmem_ram_62__15_, mem_stage_inst_dmem_ram_63__0_,
         mem_stage_inst_dmem_ram_63__1_, mem_stage_inst_dmem_ram_63__2_,
         mem_stage_inst_dmem_ram_63__3_, mem_stage_inst_dmem_ram_63__4_,
         mem_stage_inst_dmem_ram_63__5_, mem_stage_inst_dmem_ram_63__6_,
         mem_stage_inst_dmem_ram_63__7_, mem_stage_inst_dmem_ram_63__8_,
         mem_stage_inst_dmem_ram_63__9_, mem_stage_inst_dmem_ram_63__10_,
         mem_stage_inst_dmem_ram_63__11_, mem_stage_inst_dmem_ram_63__12_,
         mem_stage_inst_dmem_ram_63__13_, mem_stage_inst_dmem_ram_63__14_,
         mem_stage_inst_dmem_ram_63__15_, mem_stage_inst_dmem_ram_0__0_,
         mem_stage_inst_dmem_ram_0__1_, mem_stage_inst_dmem_ram_0__2_,
         mem_stage_inst_dmem_ram_0__3_, mem_stage_inst_dmem_ram_0__4_,
         mem_stage_inst_dmem_ram_0__5_, mem_stage_inst_dmem_ram_0__6_,
         mem_stage_inst_dmem_ram_0__7_, mem_stage_inst_dmem_ram_0__8_,
         mem_stage_inst_dmem_ram_0__9_, mem_stage_inst_dmem_ram_0__10_,
         mem_stage_inst_dmem_ram_0__11_, mem_stage_inst_dmem_ram_0__12_,
         mem_stage_inst_dmem_ram_0__13_, mem_stage_inst_dmem_ram_0__14_,
         mem_stage_inst_dmem_ram_0__15_, mem_stage_inst_dmem_ram_1__0_,
         mem_stage_inst_dmem_ram_1__1_, mem_stage_inst_dmem_ram_1__2_,
         mem_stage_inst_dmem_ram_1__3_, mem_stage_inst_dmem_ram_1__4_,
         mem_stage_inst_dmem_ram_1__5_, mem_stage_inst_dmem_ram_1__6_,
         mem_stage_inst_dmem_ram_1__7_, mem_stage_inst_dmem_ram_1__8_,
         mem_stage_inst_dmem_ram_1__9_, mem_stage_inst_dmem_ram_1__10_,
         mem_stage_inst_dmem_ram_1__11_, mem_stage_inst_dmem_ram_1__12_,
         mem_stage_inst_dmem_ram_1__13_, mem_stage_inst_dmem_ram_1__14_,
         mem_stage_inst_dmem_ram_1__15_, mem_stage_inst_dmem_ram_2__0_,
         mem_stage_inst_dmem_ram_2__1_, mem_stage_inst_dmem_ram_2__2_,
         mem_stage_inst_dmem_ram_2__3_, mem_stage_inst_dmem_ram_2__4_,
         mem_stage_inst_dmem_ram_2__5_, mem_stage_inst_dmem_ram_2__6_,
         mem_stage_inst_dmem_ram_2__7_, mem_stage_inst_dmem_ram_2__8_,
         mem_stage_inst_dmem_ram_2__9_, mem_stage_inst_dmem_ram_2__10_,
         mem_stage_inst_dmem_ram_2__11_, mem_stage_inst_dmem_ram_2__12_,
         mem_stage_inst_dmem_ram_2__13_, mem_stage_inst_dmem_ram_2__14_,
         mem_stage_inst_dmem_ram_2__15_, mem_stage_inst_dmem_ram_3__0_,
         mem_stage_inst_dmem_ram_3__1_, mem_stage_inst_dmem_ram_3__2_,
         mem_stage_inst_dmem_ram_3__3_, mem_stage_inst_dmem_ram_3__4_,
         mem_stage_inst_dmem_ram_3__5_, mem_stage_inst_dmem_ram_3__6_,
         mem_stage_inst_dmem_ram_3__7_, mem_stage_inst_dmem_ram_3__8_,
         mem_stage_inst_dmem_ram_3__9_, mem_stage_inst_dmem_ram_3__10_,
         mem_stage_inst_dmem_ram_3__11_, mem_stage_inst_dmem_ram_3__12_,
         mem_stage_inst_dmem_ram_3__13_, mem_stage_inst_dmem_ram_3__14_,
         mem_stage_inst_dmem_ram_3__15_, mem_stage_inst_dmem_ram_4__0_,
         mem_stage_inst_dmem_ram_4__1_, mem_stage_inst_dmem_ram_4__2_,
         mem_stage_inst_dmem_ram_4__3_, mem_stage_inst_dmem_ram_4__4_,
         mem_stage_inst_dmem_ram_4__5_, mem_stage_inst_dmem_ram_4__6_,
         mem_stage_inst_dmem_ram_4__7_, mem_stage_inst_dmem_ram_4__8_,
         mem_stage_inst_dmem_ram_4__9_, mem_stage_inst_dmem_ram_4__10_,
         mem_stage_inst_dmem_ram_4__11_, mem_stage_inst_dmem_ram_4__12_,
         mem_stage_inst_dmem_ram_4__13_, mem_stage_inst_dmem_ram_4__14_,
         mem_stage_inst_dmem_ram_4__15_, mem_stage_inst_dmem_ram_5__0_,
         mem_stage_inst_dmem_ram_5__1_, mem_stage_inst_dmem_ram_5__2_,
         mem_stage_inst_dmem_ram_5__3_, mem_stage_inst_dmem_ram_5__4_,
         mem_stage_inst_dmem_ram_5__5_, mem_stage_inst_dmem_ram_5__6_,
         mem_stage_inst_dmem_ram_5__7_, mem_stage_inst_dmem_ram_5__8_,
         mem_stage_inst_dmem_ram_5__9_, mem_stage_inst_dmem_ram_5__10_,
         mem_stage_inst_dmem_ram_5__11_, mem_stage_inst_dmem_ram_5__12_,
         mem_stage_inst_dmem_ram_5__13_, mem_stage_inst_dmem_ram_5__14_,
         mem_stage_inst_dmem_ram_5__15_, mem_stage_inst_dmem_ram_6__0_,
         mem_stage_inst_dmem_ram_6__1_, mem_stage_inst_dmem_ram_6__2_,
         mem_stage_inst_dmem_ram_6__3_, mem_stage_inst_dmem_ram_6__4_,
         mem_stage_inst_dmem_ram_6__5_, mem_stage_inst_dmem_ram_6__6_,
         mem_stage_inst_dmem_ram_6__7_, mem_stage_inst_dmem_ram_6__8_,
         mem_stage_inst_dmem_ram_6__9_, mem_stage_inst_dmem_ram_6__10_,
         mem_stage_inst_dmem_ram_6__11_, mem_stage_inst_dmem_ram_6__12_,
         mem_stage_inst_dmem_ram_6__13_, mem_stage_inst_dmem_ram_6__14_,
         mem_stage_inst_dmem_ram_6__15_, mem_stage_inst_dmem_ram_7__0_,
         mem_stage_inst_dmem_ram_7__1_, mem_stage_inst_dmem_ram_7__2_,
         mem_stage_inst_dmem_ram_7__3_, mem_stage_inst_dmem_ram_7__4_,
         mem_stage_inst_dmem_ram_7__5_, mem_stage_inst_dmem_ram_7__6_,
         mem_stage_inst_dmem_ram_7__7_, mem_stage_inst_dmem_ram_7__8_,
         mem_stage_inst_dmem_ram_7__9_, mem_stage_inst_dmem_ram_7__10_,
         mem_stage_inst_dmem_ram_7__11_, mem_stage_inst_dmem_ram_7__12_,
         mem_stage_inst_dmem_ram_7__13_, mem_stage_inst_dmem_ram_7__14_,
         mem_stage_inst_dmem_ram_7__15_, mem_stage_inst_dmem_ram_8__0_,
         mem_stage_inst_dmem_ram_8__1_, mem_stage_inst_dmem_ram_8__2_,
         mem_stage_inst_dmem_ram_8__3_, mem_stage_inst_dmem_ram_8__4_,
         mem_stage_inst_dmem_ram_8__5_, mem_stage_inst_dmem_ram_8__6_,
         mem_stage_inst_dmem_ram_8__7_, mem_stage_inst_dmem_ram_8__8_,
         mem_stage_inst_dmem_ram_8__9_, mem_stage_inst_dmem_ram_8__10_,
         mem_stage_inst_dmem_ram_8__11_, mem_stage_inst_dmem_ram_8__12_,
         mem_stage_inst_dmem_ram_8__13_, mem_stage_inst_dmem_ram_8__14_,
         mem_stage_inst_dmem_ram_8__15_, mem_stage_inst_dmem_ram_9__0_,
         mem_stage_inst_dmem_ram_9__1_, mem_stage_inst_dmem_ram_9__2_,
         mem_stage_inst_dmem_ram_9__3_, mem_stage_inst_dmem_ram_9__4_,
         mem_stage_inst_dmem_ram_9__5_, mem_stage_inst_dmem_ram_9__6_,
         mem_stage_inst_dmem_ram_9__7_, mem_stage_inst_dmem_ram_9__8_,
         mem_stage_inst_dmem_ram_9__9_, mem_stage_inst_dmem_ram_9__10_,
         mem_stage_inst_dmem_ram_9__11_, mem_stage_inst_dmem_ram_9__12_,
         mem_stage_inst_dmem_ram_9__13_, mem_stage_inst_dmem_ram_9__14_,
         mem_stage_inst_dmem_ram_9__15_, mem_stage_inst_dmem_ram_10__0_,
         mem_stage_inst_dmem_ram_10__1_, mem_stage_inst_dmem_ram_10__2_,
         mem_stage_inst_dmem_ram_10__3_, mem_stage_inst_dmem_ram_10__4_,
         mem_stage_inst_dmem_ram_10__5_, mem_stage_inst_dmem_ram_10__6_,
         mem_stage_inst_dmem_ram_10__7_, mem_stage_inst_dmem_ram_10__8_,
         mem_stage_inst_dmem_ram_10__9_, mem_stage_inst_dmem_ram_10__10_,
         mem_stage_inst_dmem_ram_10__11_, mem_stage_inst_dmem_ram_10__12_,
         mem_stage_inst_dmem_ram_10__13_, mem_stage_inst_dmem_ram_10__14_,
         mem_stage_inst_dmem_ram_10__15_, mem_stage_inst_dmem_ram_11__0_,
         mem_stage_inst_dmem_ram_11__1_, mem_stage_inst_dmem_ram_11__2_,
         mem_stage_inst_dmem_ram_11__3_, mem_stage_inst_dmem_ram_11__4_,
         mem_stage_inst_dmem_ram_11__5_, mem_stage_inst_dmem_ram_11__6_,
         mem_stage_inst_dmem_ram_11__7_, mem_stage_inst_dmem_ram_11__8_,
         mem_stage_inst_dmem_ram_11__9_, mem_stage_inst_dmem_ram_11__10_,
         mem_stage_inst_dmem_ram_11__11_, mem_stage_inst_dmem_ram_11__12_,
         mem_stage_inst_dmem_ram_11__13_, mem_stage_inst_dmem_ram_11__14_,
         mem_stage_inst_dmem_ram_11__15_, mem_stage_inst_dmem_ram_12__0_,
         mem_stage_inst_dmem_ram_12__1_, mem_stage_inst_dmem_ram_12__2_,
         mem_stage_inst_dmem_ram_12__3_, mem_stage_inst_dmem_ram_12__4_,
         mem_stage_inst_dmem_ram_12__5_, mem_stage_inst_dmem_ram_12__6_,
         mem_stage_inst_dmem_ram_12__7_, mem_stage_inst_dmem_ram_12__8_,
         mem_stage_inst_dmem_ram_12__9_, mem_stage_inst_dmem_ram_12__10_,
         mem_stage_inst_dmem_ram_12__11_, mem_stage_inst_dmem_ram_12__12_,
         mem_stage_inst_dmem_ram_12__13_, mem_stage_inst_dmem_ram_12__14_,
         mem_stage_inst_dmem_ram_12__15_, mem_stage_inst_dmem_ram_13__0_,
         mem_stage_inst_dmem_ram_13__1_, mem_stage_inst_dmem_ram_13__2_,
         mem_stage_inst_dmem_ram_13__3_, mem_stage_inst_dmem_ram_13__4_,
         mem_stage_inst_dmem_ram_13__5_, mem_stage_inst_dmem_ram_13__6_,
         mem_stage_inst_dmem_ram_13__7_, mem_stage_inst_dmem_ram_13__8_,
         mem_stage_inst_dmem_ram_13__9_, mem_stage_inst_dmem_ram_13__10_,
         mem_stage_inst_dmem_ram_13__11_, mem_stage_inst_dmem_ram_13__12_,
         mem_stage_inst_dmem_ram_13__13_, mem_stage_inst_dmem_ram_13__14_,
         mem_stage_inst_dmem_ram_13__15_, mem_stage_inst_dmem_ram_14__0_,
         mem_stage_inst_dmem_ram_14__1_, mem_stage_inst_dmem_ram_14__2_,
         mem_stage_inst_dmem_ram_14__3_, mem_stage_inst_dmem_ram_14__4_,
         mem_stage_inst_dmem_ram_14__5_, mem_stage_inst_dmem_ram_14__6_,
         mem_stage_inst_dmem_ram_14__7_, mem_stage_inst_dmem_ram_14__8_,
         mem_stage_inst_dmem_ram_14__9_, mem_stage_inst_dmem_ram_14__10_,
         mem_stage_inst_dmem_ram_14__11_, mem_stage_inst_dmem_ram_14__12_,
         mem_stage_inst_dmem_ram_14__13_, mem_stage_inst_dmem_ram_14__14_,
         mem_stage_inst_dmem_ram_14__15_, mem_stage_inst_dmem_ram_15__0_,
         mem_stage_inst_dmem_ram_15__1_, mem_stage_inst_dmem_ram_15__2_,
         mem_stage_inst_dmem_ram_15__3_, mem_stage_inst_dmem_ram_15__4_,
         mem_stage_inst_dmem_ram_15__5_, mem_stage_inst_dmem_ram_15__6_,
         mem_stage_inst_dmem_ram_15__7_, mem_stage_inst_dmem_ram_15__8_,
         mem_stage_inst_dmem_ram_15__9_, mem_stage_inst_dmem_ram_15__10_,
         mem_stage_inst_dmem_ram_15__11_, mem_stage_inst_dmem_ram_15__12_,
         mem_stage_inst_dmem_ram_15__13_, mem_stage_inst_dmem_ram_15__14_,
         mem_stage_inst_dmem_ram_15__15_, mem_stage_inst_dmem_ram_16__0_,
         mem_stage_inst_dmem_ram_16__1_, mem_stage_inst_dmem_ram_16__2_,
         mem_stage_inst_dmem_ram_16__3_, mem_stage_inst_dmem_ram_16__4_,
         mem_stage_inst_dmem_ram_16__5_, mem_stage_inst_dmem_ram_16__6_,
         mem_stage_inst_dmem_ram_16__7_, mem_stage_inst_dmem_ram_16__8_,
         mem_stage_inst_dmem_ram_16__9_, mem_stage_inst_dmem_ram_16__10_,
         mem_stage_inst_dmem_ram_16__11_, mem_stage_inst_dmem_ram_16__12_,
         mem_stage_inst_dmem_ram_16__13_, mem_stage_inst_dmem_ram_16__14_,
         mem_stage_inst_dmem_ram_16__15_, mem_stage_inst_dmem_ram_17__0_,
         mem_stage_inst_dmem_ram_17__1_, mem_stage_inst_dmem_ram_17__2_,
         mem_stage_inst_dmem_ram_17__3_, mem_stage_inst_dmem_ram_17__4_,
         mem_stage_inst_dmem_ram_17__5_, mem_stage_inst_dmem_ram_17__6_,
         mem_stage_inst_dmem_ram_17__7_, mem_stage_inst_dmem_ram_17__8_,
         mem_stage_inst_dmem_ram_17__9_, mem_stage_inst_dmem_ram_17__10_,
         mem_stage_inst_dmem_ram_17__11_, mem_stage_inst_dmem_ram_17__12_,
         mem_stage_inst_dmem_ram_17__13_, mem_stage_inst_dmem_ram_17__14_,
         mem_stage_inst_dmem_ram_17__15_, mem_stage_inst_dmem_ram_18__0_,
         mem_stage_inst_dmem_ram_18__1_, mem_stage_inst_dmem_ram_18__2_,
         mem_stage_inst_dmem_ram_18__3_, mem_stage_inst_dmem_ram_18__4_,
         mem_stage_inst_dmem_ram_18__5_, mem_stage_inst_dmem_ram_18__6_,
         mem_stage_inst_dmem_ram_18__7_, mem_stage_inst_dmem_ram_18__8_,
         mem_stage_inst_dmem_ram_18__9_, mem_stage_inst_dmem_ram_18__10_,
         mem_stage_inst_dmem_ram_18__11_, mem_stage_inst_dmem_ram_18__12_,
         mem_stage_inst_dmem_ram_18__13_, mem_stage_inst_dmem_ram_18__14_,
         mem_stage_inst_dmem_ram_18__15_, mem_stage_inst_dmem_ram_19__0_,
         mem_stage_inst_dmem_ram_19__1_, mem_stage_inst_dmem_ram_19__2_,
         mem_stage_inst_dmem_ram_19__3_, mem_stage_inst_dmem_ram_19__4_,
         mem_stage_inst_dmem_ram_19__5_, mem_stage_inst_dmem_ram_19__6_,
         mem_stage_inst_dmem_ram_19__7_, mem_stage_inst_dmem_ram_19__8_,
         mem_stage_inst_dmem_ram_19__9_, mem_stage_inst_dmem_ram_19__10_,
         mem_stage_inst_dmem_ram_19__11_, mem_stage_inst_dmem_ram_19__12_,
         mem_stage_inst_dmem_ram_19__13_, mem_stage_inst_dmem_ram_19__14_,
         mem_stage_inst_dmem_ram_19__15_, mem_stage_inst_dmem_ram_20__0_,
         mem_stage_inst_dmem_ram_20__1_, mem_stage_inst_dmem_ram_20__2_,
         mem_stage_inst_dmem_ram_20__3_, mem_stage_inst_dmem_ram_20__4_,
         mem_stage_inst_dmem_ram_20__5_, mem_stage_inst_dmem_ram_20__6_,
         mem_stage_inst_dmem_ram_20__7_, mem_stage_inst_dmem_ram_20__8_,
         mem_stage_inst_dmem_ram_20__9_, mem_stage_inst_dmem_ram_20__10_,
         mem_stage_inst_dmem_ram_20__11_, mem_stage_inst_dmem_ram_20__12_,
         mem_stage_inst_dmem_ram_20__13_, mem_stage_inst_dmem_ram_20__14_,
         mem_stage_inst_dmem_ram_20__15_, mem_stage_inst_dmem_ram_21__0_,
         mem_stage_inst_dmem_ram_21__1_, mem_stage_inst_dmem_ram_21__2_,
         mem_stage_inst_dmem_ram_21__3_, mem_stage_inst_dmem_ram_21__4_,
         mem_stage_inst_dmem_ram_21__5_, mem_stage_inst_dmem_ram_21__6_,
         mem_stage_inst_dmem_ram_21__7_, mem_stage_inst_dmem_ram_21__8_,
         mem_stage_inst_dmem_ram_21__9_, mem_stage_inst_dmem_ram_21__10_,
         mem_stage_inst_dmem_ram_21__11_, mem_stage_inst_dmem_ram_21__12_,
         mem_stage_inst_dmem_ram_21__13_, mem_stage_inst_dmem_ram_21__14_,
         mem_stage_inst_dmem_ram_21__15_, mem_stage_inst_dmem_ram_22__0_,
         mem_stage_inst_dmem_ram_22__1_, mem_stage_inst_dmem_ram_22__2_,
         mem_stage_inst_dmem_ram_22__3_, mem_stage_inst_dmem_ram_22__4_,
         mem_stage_inst_dmem_ram_22__5_, mem_stage_inst_dmem_ram_22__6_,
         mem_stage_inst_dmem_ram_22__7_, mem_stage_inst_dmem_ram_22__8_,
         mem_stage_inst_dmem_ram_22__9_, mem_stage_inst_dmem_ram_22__10_,
         mem_stage_inst_dmem_ram_22__11_, mem_stage_inst_dmem_ram_22__12_,
         mem_stage_inst_dmem_ram_22__13_, mem_stage_inst_dmem_ram_22__14_,
         mem_stage_inst_dmem_ram_22__15_, mem_stage_inst_dmem_ram_23__0_,
         mem_stage_inst_dmem_ram_23__1_, mem_stage_inst_dmem_ram_23__2_,
         mem_stage_inst_dmem_ram_23__3_, mem_stage_inst_dmem_ram_23__4_,
         mem_stage_inst_dmem_ram_23__5_, mem_stage_inst_dmem_ram_23__6_,
         mem_stage_inst_dmem_ram_23__7_, mem_stage_inst_dmem_ram_23__8_,
         mem_stage_inst_dmem_ram_23__9_, mem_stage_inst_dmem_ram_23__10_,
         mem_stage_inst_dmem_ram_23__11_, mem_stage_inst_dmem_ram_23__12_,
         mem_stage_inst_dmem_ram_23__13_, mem_stage_inst_dmem_ram_23__14_,
         mem_stage_inst_dmem_ram_23__15_, mem_stage_inst_dmem_ram_24__0_,
         mem_stage_inst_dmem_ram_24__1_, mem_stage_inst_dmem_ram_24__2_,
         mem_stage_inst_dmem_ram_24__3_, mem_stage_inst_dmem_ram_24__4_,
         mem_stage_inst_dmem_ram_24__5_, mem_stage_inst_dmem_ram_24__6_,
         mem_stage_inst_dmem_ram_24__7_, mem_stage_inst_dmem_ram_24__8_,
         mem_stage_inst_dmem_ram_24__9_, mem_stage_inst_dmem_ram_24__10_,
         mem_stage_inst_dmem_ram_24__11_, mem_stage_inst_dmem_ram_24__12_,
         mem_stage_inst_dmem_ram_24__13_, mem_stage_inst_dmem_ram_24__14_,
         mem_stage_inst_dmem_ram_24__15_, mem_stage_inst_dmem_ram_25__0_,
         mem_stage_inst_dmem_ram_25__1_, mem_stage_inst_dmem_ram_25__2_,
         mem_stage_inst_dmem_ram_25__3_, mem_stage_inst_dmem_ram_25__4_,
         mem_stage_inst_dmem_ram_25__5_, mem_stage_inst_dmem_ram_25__6_,
         mem_stage_inst_dmem_ram_25__7_, mem_stage_inst_dmem_ram_25__8_,
         mem_stage_inst_dmem_ram_25__9_, mem_stage_inst_dmem_ram_25__10_,
         mem_stage_inst_dmem_ram_25__11_, mem_stage_inst_dmem_ram_25__12_,
         mem_stage_inst_dmem_ram_25__13_, mem_stage_inst_dmem_ram_25__14_,
         mem_stage_inst_dmem_ram_25__15_, mem_stage_inst_dmem_ram_26__0_,
         mem_stage_inst_dmem_ram_26__1_, mem_stage_inst_dmem_ram_26__2_,
         mem_stage_inst_dmem_ram_26__3_, mem_stage_inst_dmem_ram_26__4_,
         mem_stage_inst_dmem_ram_26__5_, mem_stage_inst_dmem_ram_26__6_,
         mem_stage_inst_dmem_ram_26__7_, mem_stage_inst_dmem_ram_26__8_,
         mem_stage_inst_dmem_ram_26__9_, mem_stage_inst_dmem_ram_26__10_,
         mem_stage_inst_dmem_ram_26__11_, mem_stage_inst_dmem_ram_26__12_,
         mem_stage_inst_dmem_ram_26__13_, mem_stage_inst_dmem_ram_26__14_,
         mem_stage_inst_dmem_ram_26__15_, mem_stage_inst_dmem_ram_27__0_,
         mem_stage_inst_dmem_ram_27__1_, mem_stage_inst_dmem_ram_27__2_,
         mem_stage_inst_dmem_ram_27__3_, mem_stage_inst_dmem_ram_27__4_,
         mem_stage_inst_dmem_ram_27__5_, mem_stage_inst_dmem_ram_27__6_,
         mem_stage_inst_dmem_ram_27__7_, mem_stage_inst_dmem_ram_27__8_,
         mem_stage_inst_dmem_ram_27__9_, mem_stage_inst_dmem_ram_27__10_,
         mem_stage_inst_dmem_ram_27__11_, mem_stage_inst_dmem_ram_27__12_,
         mem_stage_inst_dmem_ram_27__13_, mem_stage_inst_dmem_ram_27__14_,
         mem_stage_inst_dmem_ram_27__15_, mem_stage_inst_dmem_ram_28__0_,
         mem_stage_inst_dmem_ram_28__1_, mem_stage_inst_dmem_ram_28__2_,
         mem_stage_inst_dmem_ram_28__3_, mem_stage_inst_dmem_ram_28__4_,
         mem_stage_inst_dmem_ram_28__5_, mem_stage_inst_dmem_ram_28__6_,
         mem_stage_inst_dmem_ram_28__7_, mem_stage_inst_dmem_ram_28__8_,
         mem_stage_inst_dmem_ram_28__9_, mem_stage_inst_dmem_ram_28__10_,
         mem_stage_inst_dmem_ram_28__11_, mem_stage_inst_dmem_ram_28__12_,
         mem_stage_inst_dmem_ram_28__13_, mem_stage_inst_dmem_ram_28__14_,
         mem_stage_inst_dmem_ram_28__15_, mem_stage_inst_dmem_ram_29__0_,
         mem_stage_inst_dmem_ram_29__1_, mem_stage_inst_dmem_ram_29__2_,
         mem_stage_inst_dmem_ram_29__3_, mem_stage_inst_dmem_ram_29__4_,
         mem_stage_inst_dmem_ram_29__5_, mem_stage_inst_dmem_ram_29__6_,
         mem_stage_inst_dmem_ram_29__7_, mem_stage_inst_dmem_ram_29__8_,
         mem_stage_inst_dmem_ram_29__9_, mem_stage_inst_dmem_ram_29__10_,
         mem_stage_inst_dmem_ram_29__11_, mem_stage_inst_dmem_ram_29__12_,
         mem_stage_inst_dmem_ram_29__13_, mem_stage_inst_dmem_ram_29__14_,
         mem_stage_inst_dmem_ram_29__15_, mem_stage_inst_dmem_ram_30__0_,
         mem_stage_inst_dmem_ram_30__1_, mem_stage_inst_dmem_ram_30__2_,
         mem_stage_inst_dmem_ram_30__3_, mem_stage_inst_dmem_ram_30__4_,
         mem_stage_inst_dmem_ram_30__5_, mem_stage_inst_dmem_ram_30__6_,
         mem_stage_inst_dmem_ram_30__7_, mem_stage_inst_dmem_ram_30__8_,
         mem_stage_inst_dmem_ram_30__9_, mem_stage_inst_dmem_ram_30__10_,
         mem_stage_inst_dmem_ram_30__11_, mem_stage_inst_dmem_ram_30__12_,
         mem_stage_inst_dmem_ram_30__13_, mem_stage_inst_dmem_ram_30__14_,
         mem_stage_inst_dmem_ram_30__15_, mem_stage_inst_dmem_ram_31__0_,
         mem_stage_inst_dmem_ram_31__1_, mem_stage_inst_dmem_ram_31__2_,
         mem_stage_inst_dmem_ram_31__3_, mem_stage_inst_dmem_ram_31__4_,
         mem_stage_inst_dmem_ram_31__5_, mem_stage_inst_dmem_ram_31__6_,
         mem_stage_inst_dmem_ram_31__7_, mem_stage_inst_dmem_ram_31__8_,
         mem_stage_inst_dmem_ram_31__9_, mem_stage_inst_dmem_ram_31__10_,
         mem_stage_inst_dmem_ram_31__11_, mem_stage_inst_dmem_ram_31__12_,
         mem_stage_inst_dmem_ram_31__13_, mem_stage_inst_dmem_ram_31__14_,
         mem_stage_inst_dmem_ram_31__15_, register_file_inst_n206,
         register_file_inst_n205, register_file_inst_n204,
         register_file_inst_n203, register_file_inst_n202,
         register_file_inst_n201, register_file_inst_n200,
         register_file_inst_n199, register_file_inst_n198,
         register_file_inst_n197, register_file_inst_n196,
         register_file_inst_n195, register_file_inst_n194,
         register_file_inst_n193, register_file_inst_n192,
         register_file_inst_n191, register_file_inst_n190,
         register_file_inst_n189, register_file_inst_n188,
         register_file_inst_n187, register_file_inst_n186,
         register_file_inst_n185, register_file_inst_n184,
         register_file_inst_n183, register_file_inst_n182,
         register_file_inst_n181, register_file_inst_n180,
         register_file_inst_n179, register_file_inst_n178,
         register_file_inst_n177, register_file_inst_n176,
         register_file_inst_n175, register_file_inst_n174,
         register_file_inst_n173, register_file_inst_n172,
         register_file_inst_n171, register_file_inst_n170,
         register_file_inst_n169, register_file_inst_n168,
         register_file_inst_n167, register_file_inst_n166,
         register_file_inst_n165, register_file_inst_n164,
         register_file_inst_n163, register_file_inst_n162,
         register_file_inst_n161, register_file_inst_n160,
         register_file_inst_n159, register_file_inst_n158,
         register_file_inst_n157, register_file_inst_n156,
         register_file_inst_n155, register_file_inst_n154,
         register_file_inst_n153, register_file_inst_n152,
         register_file_inst_n151, register_file_inst_n22,
         register_file_inst_n21, register_file_inst_n20,
         register_file_inst_n19, register_file_inst_n18,
         register_file_inst_n17, register_file_inst_n16,
         register_file_inst_n15, register_file_inst_n14,
         register_file_inst_n13, register_file_inst_n12,
         register_file_inst_n11, register_file_inst_n10, register_file_inst_n9,
         register_file_inst_n8, register_file_inst_n7, register_file_inst_n6,
         register_file_inst_n5, register_file_inst_n4, register_file_inst_n3,
         register_file_inst_n2, register_file_inst_n1, register_file_inst_n150,
         register_file_inst_n149, register_file_inst_n148,
         register_file_inst_n147, register_file_inst_n146,
         register_file_inst_n145, register_file_inst_n144,
         register_file_inst_n143, register_file_inst_n142,
         register_file_inst_n141, register_file_inst_n140,
         register_file_inst_n139, register_file_inst_n138,
         register_file_inst_n137, register_file_inst_n136,
         register_file_inst_n135, register_file_inst_n134,
         register_file_inst_n133, register_file_inst_n132,
         register_file_inst_n131, register_file_inst_n130,
         register_file_inst_n129, register_file_inst_n128,
         register_file_inst_n127, register_file_inst_n126,
         register_file_inst_n125, register_file_inst_n124,
         register_file_inst_n123, register_file_inst_n122,
         register_file_inst_n121, register_file_inst_n120,
         register_file_inst_n119, register_file_inst_n118,
         register_file_inst_n117, register_file_inst_n116,
         register_file_inst_n115, register_file_inst_n114,
         register_file_inst_n113, register_file_inst_n112,
         register_file_inst_n111, register_file_inst_n110,
         register_file_inst_n109, register_file_inst_n108,
         register_file_inst_n107, register_file_inst_n106,
         register_file_inst_n105, register_file_inst_n104,
         register_file_inst_n103, register_file_inst_n102,
         register_file_inst_n101, register_file_inst_n100,
         register_file_inst_n99, register_file_inst_n98,
         register_file_inst_n97, register_file_inst_n96,
         register_file_inst_n95, register_file_inst_n94,
         register_file_inst_n93, register_file_inst_n92,
         register_file_inst_n91, register_file_inst_n90,
         register_file_inst_n89, register_file_inst_n88,
         register_file_inst_n87, register_file_inst_n86,
         register_file_inst_n85, register_file_inst_n84,
         register_file_inst_n83, register_file_inst_n82,
         register_file_inst_n81, register_file_inst_n80,
         register_file_inst_n79, register_file_inst_n78,
         register_file_inst_n77, register_file_inst_n76,
         register_file_inst_n75, register_file_inst_n74,
         register_file_inst_n73, register_file_inst_n72,
         register_file_inst_n71, register_file_inst_n70,
         register_file_inst_n69, register_file_inst_n68,
         register_file_inst_n67, register_file_inst_n66,
         register_file_inst_n65, register_file_inst_n64,
         register_file_inst_n63, register_file_inst_n62,
         register_file_inst_n61, register_file_inst_n60,
         register_file_inst_n59, register_file_inst_n58,
         register_file_inst_n57, register_file_inst_n56,
         register_file_inst_n55, register_file_inst_n54,
         register_file_inst_n53, register_file_inst_n52,
         register_file_inst_n51, register_file_inst_n50,
         register_file_inst_n49, register_file_inst_n48,
         register_file_inst_n47, register_file_inst_n46,
         register_file_inst_n45, register_file_inst_n44,
         register_file_inst_n43, register_file_inst_n42,
         register_file_inst_n41, register_file_inst_n40,
         register_file_inst_n39, register_file_inst_n38,
         register_file_inst_n37, register_file_inst_n36,
         register_file_inst_n35, register_file_inst_n34,
         register_file_inst_n33, register_file_inst_n32,
         register_file_inst_n31, register_file_inst_n30,
         register_file_inst_n29, register_file_inst_n28,
         register_file_inst_n27, register_file_inst_n26,
         register_file_inst_n25, register_file_inst_n24,
         register_file_inst_n23, register_file_inst_n600,
         register_file_inst_n590, register_file_inst_n580,
         register_file_inst_n570, register_file_inst_n560,
         register_file_inst_n550, register_file_inst_n540,
         register_file_inst_n530, register_file_inst_n520,
         register_file_inst_n510, register_file_inst_n500,
         register_file_inst_n490, register_file_inst_n480,
         register_file_inst_n470, register_file_inst_n460,
         register_file_inst_n450, register_file_inst_n440,
         register_file_inst_n430, register_file_inst_n420,
         register_file_inst_n410, register_file_inst_n400,
         register_file_inst_n390, register_file_inst_n380,
         register_file_inst_n370, register_file_inst_n360,
         register_file_inst_n350, register_file_inst_n340,
         register_file_inst_n330, register_file_inst_n320,
         register_file_inst_n310, register_file_inst_n300,
         register_file_inst_n290, register_file_inst_reg_array_0__0_,
         register_file_inst_reg_array_0__1_,
         register_file_inst_reg_array_0__2_,
         register_file_inst_reg_array_0__3_,
         register_file_inst_reg_array_0__4_,
         register_file_inst_reg_array_0__5_,
         register_file_inst_reg_array_0__6_,
         register_file_inst_reg_array_0__7_,
         register_file_inst_reg_array_0__8_,
         register_file_inst_reg_array_0__9_,
         register_file_inst_reg_array_0__10_,
         register_file_inst_reg_array_0__11_,
         register_file_inst_reg_array_0__12_,
         register_file_inst_reg_array_0__13_,
         register_file_inst_reg_array_0__14_,
         register_file_inst_reg_array_0__15_,
         register_file_inst_reg_array_1__0_,
         register_file_inst_reg_array_1__1_,
         register_file_inst_reg_array_1__2_,
         register_file_inst_reg_array_1__3_,
         register_file_inst_reg_array_1__4_,
         register_file_inst_reg_array_1__5_,
         register_file_inst_reg_array_1__6_,
         register_file_inst_reg_array_1__7_,
         register_file_inst_reg_array_1__8_,
         register_file_inst_reg_array_1__9_,
         register_file_inst_reg_array_1__10_,
         register_file_inst_reg_array_1__11_,
         register_file_inst_reg_array_1__12_,
         register_file_inst_reg_array_1__13_,
         register_file_inst_reg_array_1__14_,
         register_file_inst_reg_array_1__15_,
         register_file_inst_reg_array_2__0_,
         register_file_inst_reg_array_2__1_,
         register_file_inst_reg_array_2__2_,
         register_file_inst_reg_array_2__3_,
         register_file_inst_reg_array_2__4_,
         register_file_inst_reg_array_2__5_,
         register_file_inst_reg_array_2__6_,
         register_file_inst_reg_array_2__7_,
         register_file_inst_reg_array_2__8_,
         register_file_inst_reg_array_2__9_,
         register_file_inst_reg_array_2__10_,
         register_file_inst_reg_array_2__11_,
         register_file_inst_reg_array_2__12_,
         register_file_inst_reg_array_2__13_,
         register_file_inst_reg_array_2__14_,
         register_file_inst_reg_array_2__15_,
         register_file_inst_reg_array_3__0_,
         register_file_inst_reg_array_3__1_,
         register_file_inst_reg_array_3__2_,
         register_file_inst_reg_array_3__3_,
         register_file_inst_reg_array_3__4_,
         register_file_inst_reg_array_3__5_,
         register_file_inst_reg_array_3__6_,
         register_file_inst_reg_array_3__7_,
         register_file_inst_reg_array_3__8_,
         register_file_inst_reg_array_3__9_,
         register_file_inst_reg_array_3__10_,
         register_file_inst_reg_array_3__11_,
         register_file_inst_reg_array_3__12_,
         register_file_inst_reg_array_3__13_,
         register_file_inst_reg_array_3__14_,
         register_file_inst_reg_array_3__15_,
         register_file_inst_reg_array_4__0_,
         register_file_inst_reg_array_4__1_,
         register_file_inst_reg_array_4__2_,
         register_file_inst_reg_array_4__3_,
         register_file_inst_reg_array_4__4_,
         register_file_inst_reg_array_4__5_,
         register_file_inst_reg_array_4__6_,
         register_file_inst_reg_array_4__7_,
         register_file_inst_reg_array_4__8_,
         register_file_inst_reg_array_4__9_,
         register_file_inst_reg_array_4__10_,
         register_file_inst_reg_array_4__11_,
         register_file_inst_reg_array_4__12_,
         register_file_inst_reg_array_4__13_,
         register_file_inst_reg_array_4__14_,
         register_file_inst_reg_array_4__15_,
         register_file_inst_reg_array_5__0_,
         register_file_inst_reg_array_5__1_,
         register_file_inst_reg_array_5__2_,
         register_file_inst_reg_array_5__3_,
         register_file_inst_reg_array_5__4_,
         register_file_inst_reg_array_5__5_,
         register_file_inst_reg_array_5__6_,
         register_file_inst_reg_array_5__7_,
         register_file_inst_reg_array_5__8_,
         register_file_inst_reg_array_5__9_,
         register_file_inst_reg_array_5__10_,
         register_file_inst_reg_array_5__11_,
         register_file_inst_reg_array_5__12_,
         register_file_inst_reg_array_5__13_,
         register_file_inst_reg_array_5__14_,
         register_file_inst_reg_array_5__15_,
         register_file_inst_reg_array_6__0_,
         register_file_inst_reg_array_6__1_,
         register_file_inst_reg_array_6__2_,
         register_file_inst_reg_array_6__3_,
         register_file_inst_reg_array_6__4_,
         register_file_inst_reg_array_6__5_,
         register_file_inst_reg_array_6__6_,
         register_file_inst_reg_array_6__7_,
         register_file_inst_reg_array_6__8_,
         register_file_inst_reg_array_6__9_,
         register_file_inst_reg_array_6__10_,
         register_file_inst_reg_array_6__11_,
         register_file_inst_reg_array_6__12_,
         register_file_inst_reg_array_6__13_,
         register_file_inst_reg_array_6__14_,
         register_file_inst_reg_array_6__15_,
         register_file_inst_reg_array_7__0_,
         register_file_inst_reg_array_7__1_,
         register_file_inst_reg_array_7__2_,
         register_file_inst_reg_array_7__3_,
         register_file_inst_reg_array_7__4_,
         register_file_inst_reg_array_7__5_,
         register_file_inst_reg_array_7__6_,
         register_file_inst_reg_array_7__7_,
         register_file_inst_reg_array_7__8_,
         register_file_inst_reg_array_7__9_,
         register_file_inst_reg_array_7__10_,
         register_file_inst_reg_array_7__11_,
         register_file_inst_reg_array_7__12_,
         register_file_inst_reg_array_7__13_,
         register_file_inst_reg_array_7__14_,
         register_file_inst_reg_array_7__15_, hazard_detection_unit_inst_n32,
         hazard_detection_unit_inst_n31, hazard_detection_unit_inst_n30,
         hazard_detection_unit_inst_n29, hazard_detection_unit_inst_n28,
         hazard_detection_unit_inst_n27, hazard_detection_unit_inst_n26,
         hazard_detection_unit_inst_n25, hazard_detection_unit_inst_n24,
         hazard_detection_unit_inst_n23, hazard_detection_unit_inst_n22,
         hazard_detection_unit_inst_n21, hazard_detection_unit_inst_n20,
         hazard_detection_unit_inst_n19, hazard_detection_unit_inst_n18,
         hazard_detection_unit_inst_n17, hazard_detection_unit_inst_n16,
         hazard_detection_unit_inst_n15, hazard_detection_unit_inst_n14,
         hazard_detection_unit_inst_n13, hazard_detection_unit_inst_n12,
         hazard_detection_unit_inst_n11, hazard_detection_unit_inst_n10,
         hazard_detection_unit_inst_n9, hazard_detection_unit_inst_n8,
         hazard_detection_unit_inst_n7, hazard_detection_unit_inst_n6,
         hazard_detection_unit_inst_n5, hazard_detection_unit_inst_n4,
         hazard_detection_unit_inst_n3, hazard_detection_unit_inst_n2,
         hazard_detection_unit_inst_n1;
  wire   [5:0] branch_offset_imm;
  wire   [56:0] id_pipeline_reg_out;
  wire   [2:0] reg_read_addr_1;
  wire   [2:0] reg_read_addr_2;
  wire   [15:0] reg_read_data_1;
  wire   [15:0] reg_read_data_2;
  wire   [2:0] decoding_op_src2;
  wire   [37:0] ex_pipeline_reg_out;
  wire   [2:0] ex_op_dest;
  wire   [36:0] mem_pipeline_reg_out;
  wire   [2:0] mem_op_dest;
  wire   [2:0] reg_write_dest;
  wire   [15:0] reg_write_data;
  wire   [7:2] if_stage_inst_r301_carry;
  wire   [15:0] id_stage_inst_ex_alu_src2;
  wire   [2:0] id_stage_inst_ex_alu_cmd;
  wire   [15:0] ex_stage_inst_ex_alu_result;
  wire   [15:0] ex_stage_inst_alu_inst_r316_b_as;
  wire   [15:0] mem_stage_inst_mem_read_data;
  wire   rst;

  TIELO_X1M_A12TS rst_node ( .Y(rst) );
  TIELO_X1M_A12TS u1 ( .Y(n1) );
  NAND2B_X0P5M_A12TS if_stage_inst_u17 ( .AN(branch_offset_imm[0]), .B(
        branch_taken), .Y(if_stage_inst_u3_u1_z_0) );
  AND2_X0P5M_A12TS if_stage_inst_u16 ( .A(branch_offset_imm[1]), .B(
        branch_taken), .Y(if_stage_inst_u3_u1_z_1) );
  AND2_X0P5M_A12TS if_stage_inst_u15 ( .A(branch_offset_imm[2]), .B(
        branch_taken), .Y(if_stage_inst_u3_u1_z_2) );
  AND2_X0P5M_A12TS if_stage_inst_u14 ( .A(branch_offset_imm[3]), .B(
        branch_taken), .Y(if_stage_inst_u3_u1_z_3) );
  AND2_X0P5M_A12TS if_stage_inst_u13 ( .A(branch_offset_imm[4]), .B(
        branch_taken), .Y(if_stage_inst_u3_u1_z_4) );
  AND2_X0P5M_A12TS if_stage_inst_u12 ( .A(branch_taken), .B(
        branch_offset_imm[5]), .Y(if_stage_inst_u3_u1_z_7) );
  MXT2_X0P5M_A12TS if_stage_inst_u11 ( .A(pc[7]), .B(if_stage_inst_n29), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n12) );
  MXT2_X0P5M_A12TS if_stage_inst_u10 ( .A(pc[6]), .B(if_stage_inst_n28), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n13) );
  MXT2_X0P5M_A12TS if_stage_inst_u9 ( .A(pc[5]), .B(if_stage_inst_n27), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n14) );
  MXT2_X0P5M_A12TS if_stage_inst_u8 ( .A(pc[4]), .B(if_stage_inst_n26), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n15) );
  MXT2_X0P5M_A12TS if_stage_inst_u7 ( .A(pc[3]), .B(if_stage_inst_n25), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n16) );
  MXT2_X0P5M_A12TS if_stage_inst_u6 ( .A(pc[2]), .B(if_stage_inst_n24), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n17) );
  MXT2_X0P5M_A12TS if_stage_inst_u5 ( .A(pc[1]), .B(if_stage_inst_n23), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n18) );
  MXT2_X0P5M_A12TS if_stage_inst_u4 ( .A(pc[0]), .B(if_stage_inst_n22), .S0(
        pipeline_stall_n), .Y(if_stage_inst_n19) );
  TIELO_X1M_A12TS if_stage_inst_u3 ( .Y(if_stage_inst_instruction_0_) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_0_ ( .D(if_stage_inst_n19), .CK(clk), 
        .R(rst), .Q(pc[0]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_7_ ( .D(if_stage_inst_n12), .CK(clk), 
        .R(rst), .Q(pc[7]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_6_ ( .D(if_stage_inst_n13), .CK(clk), 
        .R(rst), .Q(pc[6]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_5_ ( .D(if_stage_inst_n14), .CK(clk), 
        .R(rst), .Q(pc[5]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_4_ ( .D(if_stage_inst_n15), .CK(clk), 
        .R(rst), .Q(pc[4]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_3_ ( .D(if_stage_inst_n16), .CK(clk), 
        .R(rst), .Q(pc[3]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_2_ ( .D(if_stage_inst_n17), .CK(clk), 
        .R(rst), .Q(pc[2]) );
  DFFRPQ_X1M_A12TS if_stage_inst_pc_reg_1_ ( .D(if_stage_inst_n18), .CK(clk), 
        .R(rst), .Q(pc[1]) );
  TIELO_X1M_A12TS if_stage_inst_imem_u2 ( .Y(
        if_stage_inst_imem_instruction_15_) );
  AND2_X1M_A12TS if_stage_inst_r301_u2 ( .A(if_stage_inst_u3_u1_z_0), .B(pc[0]), .Y(if_stage_inst_r301_n1) );
  XOR2_X1M_A12TS if_stage_inst_r301_u1 ( .A(if_stage_inst_u3_u1_z_0), .B(pc[0]), .Y(if_stage_inst_n22) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_1 ( .A(pc[1]), .B(
        if_stage_inst_u3_u1_z_1), .CI(if_stage_inst_r301_n1), .CO(
        if_stage_inst_r301_carry[2]), .S(if_stage_inst_n23) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_2 ( .A(pc[2]), .B(
        if_stage_inst_u3_u1_z_2), .CI(if_stage_inst_r301_carry[2]), .CO(
        if_stage_inst_r301_carry[3]), .S(if_stage_inst_n24) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_3 ( .A(pc[3]), .B(
        if_stage_inst_u3_u1_z_3), .CI(if_stage_inst_r301_carry[3]), .CO(
        if_stage_inst_r301_carry[4]), .S(if_stage_inst_n25) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_4 ( .A(pc[4]), .B(
        if_stage_inst_u3_u1_z_4), .CI(if_stage_inst_r301_carry[4]), .CO(
        if_stage_inst_r301_carry[5]), .S(if_stage_inst_n26) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_5 ( .A(pc[5]), .B(
        if_stage_inst_u3_u1_z_7), .CI(if_stage_inst_r301_carry[5]), .CO(
        if_stage_inst_r301_carry[6]), .S(if_stage_inst_n27) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_6 ( .A(pc[6]), .B(
        if_stage_inst_u3_u1_z_7), .CI(if_stage_inst_r301_carry[6]), .CO(
        if_stage_inst_r301_carry[7]), .S(if_stage_inst_n28) );
  ADDF_X1M_A12TS if_stage_inst_r301_u1_7 ( .A(pc[7]), .B(
        if_stage_inst_u3_u1_z_7), .CI(if_stage_inst_r301_carry[7]), .CO(), .S(
        if_stage_inst_n29) );
  OR6_X0P5M_A12TS id_stage_inst_u92 ( .A(reg_read_data_1[6]), .B(
        reg_read_data_1[5]), .C(reg_read_data_1[4]), .D(reg_read_data_1[9]), 
        .E(reg_read_data_1[8]), .F(reg_read_data_1[7]), .Y(id_stage_inst_n42)
         );
  OR6_X0P5M_A12TS id_stage_inst_u91 ( .A(reg_read_data_1[3]), .B(
        reg_read_data_1[2]), .C(reg_read_data_1[1]), .D(reg_read_data_1[15]), 
        .E(reg_read_data_1[14]), .F(id_stage_inst_n42), .Y(id_stage_inst_n38)
         );
  OR6_X0P5M_A12TS id_stage_inst_u90 ( .A(reg_read_data_1[10]), .B(
        reg_read_data_1[0]), .C(id_stage_inst_n44), .D(reg_read_data_1[13]), 
        .E(reg_read_data_1[12]), .F(reg_read_data_1[11]), .Y(id_stage_inst_n39) );
  NAND2_X0P5A_A12TS id_stage_inst_u89 ( .A(id_stage_inst_instruction_reg_10_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n9) );
  NAND2_X0P5A_A12TS id_stage_inst_u88 ( .A(id_stage_inst_instruction_reg_11_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n8) );
  INV_X0P5B_A12TS id_stage_inst_u87 ( .A(id_stage_inst_instruction_reg_14_), 
        .Y(id_stage_inst_n37) );
  OR2_X0P5M_A12TS id_stage_inst_u86 ( .A(id_stage_inst_instruction_reg_13_), 
        .B(id_stage_inst_instruction_reg_12_), .Y(id_stage_inst_n36) );
  NOR2_X0P5A_A12TS id_stage_inst_u85 ( .A(id_stage_inst_n37), .B(
        id_stage_inst_n36), .Y(id_stage_inst_n41) );
  NAND4_X0P5A_A12TS id_stage_inst_u84 ( .A(id_stage_inst_n9), .B(
        id_stage_inst_n8), .C(id_stage_inst_instruction_reg_15_), .D(
        id_stage_inst_n41), .Y(id_stage_inst_n40) );
  NOR3_X0P5A_A12TS id_stage_inst_u83 ( .A(id_stage_inst_n38), .B(
        id_stage_inst_n39), .C(id_stage_inst_n40), .Y(branch_taken) );
  AND4_X0P5M_A12TS id_stage_inst_u82 ( .A(id_stage_inst_instruction_reg_12_), 
        .B(id_stage_inst_instruction_reg_15_), .C(
        id_stage_inst_instruction_reg_13_), .D(id_stage_inst_n37), .Y(
        id_stage_inst_n66) );
  MXIT2_X0P5M_A12TS id_stage_inst_u81 ( .A(branch_offset_imm[3]), .B(
        id_stage_inst_instruction_reg_9_), .S0(id_stage_inst_n66), .Y(
        id_stage_inst_n10) );
  NOR2_X0P5A_A12TS id_stage_inst_u80 ( .A(id_stage_inst_instruction_reg_14_), 
        .B(id_stage_inst_n36), .Y(id_stage_inst_n33) );
  XNOR2_X0P5M_A12TS id_stage_inst_u79 ( .A(id_stage_inst_instruction_reg_12_), 
        .B(id_stage_inst_instruction_reg_13_), .Y(id_stage_inst_n35) );
  MXIT2_X0P5M_A12TS id_stage_inst_u78 ( .A(id_stage_inst_n35), .B(
        id_stage_inst_n36), .S0(id_stage_inst_instruction_reg_14_), .Y(
        id_stage_inst_n34) );
  MXT2_X0P5M_A12TS id_stage_inst_u77 ( .A(id_stage_inst_n33), .B(
        id_stage_inst_n34), .S0(id_stage_inst_instruction_reg_15_), .Y(
        id_stage_inst_n32) );
  NOR2_X0P5A_A12TS id_stage_inst_u76 ( .A(id_stage_inst_n10), .B(
        id_stage_inst_n32), .Y(decoding_op_src2[0]) );
  MXIT2_X0P5M_A12TS id_stage_inst_u75 ( .A(branch_offset_imm[4]), .B(
        id_stage_inst_instruction_reg_10_), .S0(id_stage_inst_n66), .Y(
        id_stage_inst_n11) );
  NOR2_X0P5A_A12TS id_stage_inst_u74 ( .A(id_stage_inst_n11), .B(
        id_stage_inst_n32), .Y(decoding_op_src2[1]) );
  MXIT2_X0P5M_A12TS id_stage_inst_u73 ( .A(branch_offset_imm[5]), .B(
        id_stage_inst_instruction_reg_11_), .S0(id_stage_inst_n66), .Y(
        id_stage_inst_n12) );
  NOR2_X0P5A_A12TS id_stage_inst_u72 ( .A(id_stage_inst_n12), .B(
        id_stage_inst_n32), .Y(decoding_op_src2[2]) );
  NAND2_X0P5A_A12TS id_stage_inst_u71 ( .A(id_stage_inst_instruction_reg_15_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n2) );
  INV_X0P5B_A12TS id_stage_inst_u70 ( .A(rst), .Y(id_stage_inst_n6) );
  NAND2_X0P5A_A12TS id_stage_inst_u69 ( .A(id_stage_inst_n2), .B(
        id_stage_inst_n6), .Y(id_stage_inst_n28) );
  NAND2_X0P5A_A12TS id_stage_inst_u68 ( .A(id_stage_inst_instruction_reg_12_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n17) );
  INV_X0P5B_A12TS id_stage_inst_u67 ( .A(id_stage_inst_n17), .Y(
        id_stage_inst_n24) );
  NAND2_X0P5A_A12TS id_stage_inst_u66 ( .A(id_stage_inst_instruction_reg_13_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n26) );
  INV_X0P5B_A12TS id_stage_inst_u65 ( .A(id_stage_inst_n26), .Y(
        id_stage_inst_n31) );
  NAND2_X0P5A_A12TS id_stage_inst_u64 ( .A(id_stage_inst_instruction_reg_14_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n27) );
  INV_X0P5B_A12TS id_stage_inst_u63 ( .A(id_stage_inst_n27), .Y(
        id_stage_inst_n25) );
  NOR2_X0P5A_A12TS id_stage_inst_u62 ( .A(id_stage_inst_n31), .B(
        id_stage_inst_n25), .Y(id_stage_inst_n22) );
  INV_X0P5B_A12TS id_stage_inst_u61 ( .A(id_stage_inst_n2), .Y(
        id_stage_inst_n23) );
  NOR2_X0P5A_A12TS id_stage_inst_u60 ( .A(id_stage_inst_n24), .B(
        id_stage_inst_n31), .Y(id_stage_inst_n19) );
  NOR2B_X0P5M_A12TS id_stage_inst_u59 ( .AN(id_stage_inst_n19), .B(
        id_stage_inst_n25), .Y(id_stage_inst_n1) );
  NAND3_X0P5A_A12TS id_stage_inst_u58 ( .A(id_stage_inst_n23), .B(
        id_stage_inst_n6), .C(id_stage_inst_n1), .Y(id_stage_inst_n29) );
  OAI31_X0P5M_A12TS id_stage_inst_u57 ( .A0(id_stage_inst_n28), .A1(
        id_stage_inst_n24), .A2(id_stage_inst_n22), .B0(id_stage_inst_n29), 
        .Y(id_stage_inst_ex_alu_cmd[0]) );
  AOI22_X0P5M_A12TS id_stage_inst_u56 ( .A0(id_stage_inst_n19), .A1(
        id_stage_inst_n25), .B0(id_stage_inst_n24), .B1(id_stage_inst_n31), 
        .Y(id_stage_inst_n30) );
  OAI21_X0P5M_A12TS id_stage_inst_u55 ( .A0(id_stage_inst_n30), .A1(
        id_stage_inst_n28), .B0(id_stage_inst_n29), .Y(
        id_stage_inst_ex_alu_cmd[1]) );
  OAI31_X0P5M_A12TS id_stage_inst_u54 ( .A0(id_stage_inst_n28), .A1(
        id_stage_inst_n19), .A2(id_stage_inst_n27), .B0(id_stage_inst_n29), 
        .Y(id_stage_inst_ex_alu_cmd[2]) );
  NOR2_X0P5A_A12TS id_stage_inst_u53 ( .A(id_stage_inst_n27), .B(
        id_stage_inst_n2), .Y(id_stage_inst_n4) );
  NOR3_X0P5A_A12TS id_stage_inst_u52 ( .A(id_stage_inst_n2), .B(
        id_stage_inst_n25), .C(id_stage_inst_n26), .Y(id_stage_inst_n18) );
  NAND2_X0P5A_A12TS id_stage_inst_u51 ( .A(id_stage_inst_n18), .B(
        id_stage_inst_n24), .Y(id_stage_inst_n5) );
  INV_X0P5B_A12TS id_stage_inst_u50 ( .A(id_stage_inst_n5), .Y(
        id_stage_inst_n20) );
  AND3_X0P5M_A12TS id_stage_inst_u49 ( .A(id_stage_inst_n22), .B(
        id_stage_inst_n23), .C(id_stage_inst_n24), .Y(id_stage_inst_n21) );
  AOI211_X0P5M_A12TS id_stage_inst_u48 ( .A0(id_stage_inst_n4), .A1(
        id_stage_inst_n19), .B0(id_stage_inst_n20), .C0(id_stage_inst_n21), 
        .Y(id_stage_inst_n16) );
  NAND3_X0P5A_A12TS id_stage_inst_u47 ( .A(id_stage_inst_n17), .B(
        id_stage_inst_n6), .C(id_stage_inst_n18), .Y(id_stage_inst_n7) );
  OAI21_X0P5M_A12TS id_stage_inst_u46 ( .A0(rst), .A1(id_stage_inst_n16), .B0(
        id_stage_inst_n7), .Y(id_stage_inst_n15) );
  INV_X0P5B_A12TS id_stage_inst_u45 ( .A(id_stage_inst_n15), .Y(
        id_stage_inst_n13) );
  MXT2_X0P5M_A12TS id_stage_inst_u44 ( .A(branch_offset_imm[0]), .B(
        reg_read_data_2[0]), .S0(id_stage_inst_n13), .Y(
        id_stage_inst_ex_alu_src2[0]) );
  NAND2_X0P5A_A12TS id_stage_inst_u43 ( .A(branch_offset_imm[5]), .B(
        id_stage_inst_n15), .Y(id_stage_inst_n14) );
  AO1B2_X0P5M_A12TS id_stage_inst_u42 ( .B0(reg_read_data_2[10]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[10]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u41 ( .B0(reg_read_data_2[11]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[11]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u40 ( .B0(reg_read_data_2[12]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[12]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u39 ( .B0(reg_read_data_2[13]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[13]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u38 ( .B0(reg_read_data_2[14]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[14]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u37 ( .B0(reg_read_data_2[15]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[15]) );
  MXT2_X0P5M_A12TS id_stage_inst_u36 ( .A(branch_offset_imm[1]), .B(
        reg_read_data_2[1]), .S0(id_stage_inst_n13), .Y(
        id_stage_inst_ex_alu_src2[1]) );
  MXT2_X0P5M_A12TS id_stage_inst_u35 ( .A(branch_offset_imm[2]), .B(
        reg_read_data_2[2]), .S0(id_stage_inst_n13), .Y(
        id_stage_inst_ex_alu_src2[2]) );
  MXT2_X0P5M_A12TS id_stage_inst_u34 ( .A(branch_offset_imm[3]), .B(
        reg_read_data_2[3]), .S0(id_stage_inst_n13), .Y(
        id_stage_inst_ex_alu_src2[3]) );
  MXT2_X0P5M_A12TS id_stage_inst_u33 ( .A(branch_offset_imm[4]), .B(
        reg_read_data_2[4]), .S0(id_stage_inst_n13), .Y(
        id_stage_inst_ex_alu_src2[4]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u32 ( .B0(reg_read_data_2[5]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[5]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u31 ( .B0(reg_read_data_2[6]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[6]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u30 ( .B0(reg_read_data_2[7]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[7]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u29 ( .B0(reg_read_data_2[8]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[8]) );
  AO1B2_X0P5M_A12TS id_stage_inst_u28 ( .B0(reg_read_data_2[9]), .B1(
        id_stage_inst_n13), .A0N(id_stage_inst_n14), .Y(
        id_stage_inst_ex_alu_src2[9]) );
  MXT2_X0P5M_A12TS id_stage_inst_u27 ( .A(branch_offset_imm[0]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n49) );
  MXT2_X0P5M_A12TS id_stage_inst_u26 ( .A(branch_offset_imm[1]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n50) );
  MXT2_X0P5M_A12TS id_stage_inst_u25 ( .A(branch_offset_imm[2]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n51) );
  MXT2_X0P5M_A12TS id_stage_inst_u24 ( .A(branch_offset_imm[3]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n52) );
  MXT2_X0P5M_A12TS id_stage_inst_u23 ( .A(branch_offset_imm[4]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n53) );
  MXT2_X0P5M_A12TS id_stage_inst_u22 ( .A(branch_offset_imm[5]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n54) );
  MXT2_X0P5M_A12TS id_stage_inst_u21 ( .A(reg_read_addr_1[0]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n55) );
  MXT2_X0P5M_A12TS id_stage_inst_u20 ( .A(reg_read_addr_1[1]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n56) );
  MXT2_X0P5M_A12TS id_stage_inst_u19 ( .A(reg_read_addr_1[2]), .B(n1), .S0(
        pipeline_stall_n), .Y(id_stage_inst_n57) );
  MXT2_X0P5M_A12TS id_stage_inst_u18 ( .A(id_stage_inst_instruction_reg_9_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n58) );
  MXT2_X0P5M_A12TS id_stage_inst_u17 ( .A(id_stage_inst_instruction_reg_10_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n59) );
  MXT2_X0P5M_A12TS id_stage_inst_u16 ( .A(id_stage_inst_instruction_reg_11_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n60) );
  MXT2_X0P5M_A12TS id_stage_inst_u15 ( .A(id_stage_inst_instruction_reg_12_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n61) );
  MXT2_X0P5M_A12TS id_stage_inst_u14 ( .A(id_stage_inst_instruction_reg_13_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n62) );
  MXT2_X0P5M_A12TS id_stage_inst_u13 ( .A(id_stage_inst_instruction_reg_14_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n63) );
  MXT2_X0P5M_A12TS id_stage_inst_u12 ( .A(id_stage_inst_instruction_reg_15_), 
        .B(n1), .S0(pipeline_stall_n), .Y(id_stage_inst_n64) );
  INV_X0P5B_A12TS id_stage_inst_u11 ( .A(id_stage_inst_n12), .Y(
        reg_read_addr_2[2]) );
  INV_X0P5B_A12TS id_stage_inst_u10 ( .A(id_stage_inst_n9), .Y(
        id_stage_inst_n46) );
  INV_X0P5B_A12TS id_stage_inst_u9 ( .A(id_stage_inst_n8), .Y(
        id_stage_inst_n45) );
  INV_X0P5B_A12TS id_stage_inst_u8 ( .A(id_stage_inst_n7), .Y(
        id_stage_inst_n43) );
  NAND2_X0P5A_A12TS id_stage_inst_u7 ( .A(id_stage_inst_n5), .B(
        id_stage_inst_n6), .Y(id_stage_inst_n3) );
  AOI211_X0P5M_A12TS id_stage_inst_u6 ( .A0(id_stage_inst_n1), .A1(
        id_stage_inst_n2), .B0(id_stage_inst_n3), .C0(id_stage_inst_n4), .Y(
        id_stage_inst_write_back_en) );
  AND2_X0P7M_A12TS id_stage_inst_u5 ( .A(id_stage_inst_instruction_reg_9_), 
        .B(pipeline_stall_n), .Y(id_stage_inst_n44) );
  INV_X1M_A12TS id_stage_inst_u4 ( .A(id_stage_inst_n10), .Y(
        reg_read_addr_2[0]) );
  INV_X1M_A12TS id_stage_inst_u3 ( .A(id_stage_inst_n11), .Y(
        reg_read_addr_2[1]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_25_ ( .D(
        id_stage_inst_ex_alu_src2[3]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[25]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_23_ ( .D(
        id_stage_inst_ex_alu_src2[1]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[23]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_22_ ( .D(
        id_stage_inst_ex_alu_src2[0]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[22]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_24_ ( .D(
        id_stage_inst_ex_alu_src2[2]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[24]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_26_ ( .D(
        id_stage_inst_ex_alu_src2[4]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[26]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_8_ ( .D(id_stage_inst_n57), .CK(clk), .R(rst), .Q(reg_read_addr_1[2]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_7_ ( .D(id_stage_inst_n56), .CK(clk), .R(rst), .Q(reg_read_addr_1[1]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_6_ ( .D(id_stage_inst_n55), .CK(clk), .R(rst), .Q(reg_read_addr_1[0]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_53_ ( .D(
        reg_read_data_1[15]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[53])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_48_ ( .D(
        reg_read_data_1[10]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[48])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_47_ ( .D(
        reg_read_data_1[9]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[47]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_49_ ( .D(
        reg_read_data_1[11]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[49])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_44_ ( .D(
        reg_read_data_1[6]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[44]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_52_ ( .D(
        reg_read_data_1[14]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[52])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_51_ ( .D(
        reg_read_data_1[13]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[51])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_40_ ( .D(
        reg_read_data_1[2]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[40]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_41_ ( .D(
        reg_read_data_1[3]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[41]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_42_ ( .D(
        reg_read_data_1[4]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[42]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_45_ ( .D(
        reg_read_data_1[7]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[45]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_43_ ( .D(
        reg_read_data_1[5]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[43]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_46_ ( .D(
        reg_read_data_1[8]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[46]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_39_ ( .D(
        reg_read_data_1[1]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[39]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_50_ ( .D(
        reg_read_data_1[12]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[50])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_38_ ( .D(
        reg_read_data_1[0]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[38]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_37_ ( .D(
        id_stage_inst_ex_alu_src2[15]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[37]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_54_ ( .D(
        id_stage_inst_ex_alu_cmd[0]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[54]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_31_ ( .D(
        id_stage_inst_ex_alu_src2[9]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[31]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_29_ ( .D(
        id_stage_inst_ex_alu_src2[7]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[29]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_27_ ( .D(
        id_stage_inst_ex_alu_src2[5]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[27]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_28_ ( .D(
        id_stage_inst_ex_alu_src2[6]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[28]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_30_ ( .D(
        id_stage_inst_ex_alu_src2[8]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[30]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_36_ ( .D(
        id_stage_inst_ex_alu_src2[14]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[36]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_35_ ( .D(
        id_stage_inst_ex_alu_src2[13]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[35]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_33_ ( .D(
        id_stage_inst_ex_alu_src2[11]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[33]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_34_ ( .D(
        id_stage_inst_ex_alu_src2[12]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[34]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_32_ ( .D(
        id_stage_inst_ex_alu_src2[10]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[32]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_14_ ( .D(
        id_stage_inst_n63), .CK(clk), .R(rst), .Q(
        id_stage_inst_instruction_reg_14_) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_12_ ( .D(
        id_stage_inst_n61), .CK(clk), .R(rst), .Q(
        id_stage_inst_instruction_reg_12_) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_15_ ( .D(
        id_stage_inst_n64), .CK(clk), .R(rst), .Q(
        id_stage_inst_instruction_reg_15_) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_13_ ( .D(
        id_stage_inst_n62), .CK(clk), .R(rst), .Q(
        id_stage_inst_instruction_reg_13_) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_1_ ( .D(
        id_stage_inst_n44), .CK(clk), .R(rst), .Q(ex_op_dest[0]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_2_ ( .D(
        id_stage_inst_n46), .CK(clk), .R(rst), .Q(ex_op_dest[1]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_3_ ( .D(
        id_stage_inst_n45), .CK(clk), .R(rst), .Q(ex_op_dest[2]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_55_ ( .D(
        id_stage_inst_ex_alu_cmd[1]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[55]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_5_ ( .D(id_stage_inst_n54), .CK(clk), .R(rst), .Q(branch_offset_imm[5]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_3_ ( .D(id_stage_inst_n52), .CK(clk), .R(rst), .Q(branch_offset_imm[3]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_4_ ( .D(id_stage_inst_n53), .CK(clk), .R(rst), .Q(branch_offset_imm[4]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_56_ ( .D(
        id_stage_inst_ex_alu_cmd[2]), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[56]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_10_ ( .D(
        id_stage_inst_n59), .CK(clk), .R(rst), .Q(
        id_stage_inst_instruction_reg_10_) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_11_ ( .D(
        id_stage_inst_n60), .CK(clk), .R(rst), .Q(
        id_stage_inst_instruction_reg_11_) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_9_ ( .D(id_stage_inst_n58), .CK(clk), .R(rst), .Q(id_stage_inst_instruction_reg_9_) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_0_ ( .D(id_stage_inst_n49), .CK(clk), .R(rst), .Q(branch_offset_imm[0]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_1_ ( .D(id_stage_inst_n50), .CK(clk), .R(rst), .Q(branch_offset_imm[1]) );
  DFFRPQ_X1M_A12TS id_stage_inst_instruction_reg_reg_2_ ( .D(id_stage_inst_n51), .CK(clk), .R(rst), .Q(branch_offset_imm[2]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_0_ ( .D(
        id_stage_inst_n43), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[0]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_4_ ( .D(
        id_stage_inst_write_back_en), .CK(clk), .R(rst), .Q(
        id_pipeline_reg_out[4]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_5_ ( .D(
        reg_read_data_2[0]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[5]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_6_ ( .D(
        reg_read_data_2[1]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[6]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_7_ ( .D(
        reg_read_data_2[2]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[7]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_8_ ( .D(
        reg_read_data_2[3]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[8]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_9_ ( .D(
        reg_read_data_2[4]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[9]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_10_ ( .D(
        reg_read_data_2[5]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[10]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_11_ ( .D(
        reg_read_data_2[6]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[11]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_12_ ( .D(
        reg_read_data_2[7]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[12]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_13_ ( .D(
        reg_read_data_2[8]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[13]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_14_ ( .D(
        reg_read_data_2[9]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[14]) );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_15_ ( .D(
        reg_read_data_2[10]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[15])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_16_ ( .D(
        reg_read_data_2[11]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[16])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_17_ ( .D(
        reg_read_data_2[12]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[17])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_18_ ( .D(
        reg_read_data_2[13]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[18])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_19_ ( .D(
        reg_read_data_2[14]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[19])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_20_ ( .D(
        reg_read_data_2[15]), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[20])
         );
  DFFRPQ_X1M_A12TS id_stage_inst_pipeline_reg_out_reg_21_ ( .D(
        id_stage_inst_n66), .CK(clk), .R(rst), .Q(id_pipeline_reg_out[21]) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u40 ( .AN(id_pipeline_reg_out[7]), .B(rst), 
        .Y(ex_stage_inst_n10) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u39 ( .AN(id_pipeline_reg_out[8]), .B(rst), 
        .Y(ex_stage_inst_n11) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u38 ( .AN(id_pipeline_reg_out[9]), .B(rst), 
        .Y(ex_stage_inst_n12) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u37 ( .AN(id_pipeline_reg_out[10]), .B(rst), 
        .Y(ex_stage_inst_n13) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u36 ( .AN(id_pipeline_reg_out[11]), .B(rst), 
        .Y(ex_stage_inst_n14) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u35 ( .AN(id_pipeline_reg_out[12]), .B(rst), 
        .Y(ex_stage_inst_n15) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u34 ( .AN(id_pipeline_reg_out[13]), .B(rst), 
        .Y(ex_stage_inst_n16) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u33 ( .AN(id_pipeline_reg_out[14]), .B(rst), 
        .Y(ex_stage_inst_n17) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u32 ( .AN(id_pipeline_reg_out[15]), .B(rst), 
        .Y(ex_stage_inst_n18) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u31 ( .AN(id_pipeline_reg_out[16]), .B(rst), 
        .Y(ex_stage_inst_n19) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u30 ( .AN(id_pipeline_reg_out[17]), .B(rst), 
        .Y(ex_stage_inst_n20) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u29 ( .AN(id_pipeline_reg_out[18]), .B(rst), 
        .Y(ex_stage_inst_n21) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u28 ( .AN(id_pipeline_reg_out[19]), .B(rst), 
        .Y(ex_stage_inst_n22) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u27 ( .AN(id_pipeline_reg_out[20]), .B(rst), 
        .Y(ex_stage_inst_n23) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u26 ( .AN(id_pipeline_reg_out[21]), .B(rst), 
        .Y(ex_stage_inst_n24) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u25 ( .AN(ex_stage_inst_ex_alu_result[0]), 
        .B(rst), .Y(ex_stage_inst_n25) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u24 ( .AN(ex_stage_inst_ex_alu_result[1]), 
        .B(rst), .Y(ex_stage_inst_n26) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u23 ( .AN(ex_stage_inst_ex_alu_result[2]), 
        .B(rst), .Y(ex_stage_inst_n27) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u22 ( .AN(ex_stage_inst_ex_alu_result[3]), 
        .B(rst), .Y(ex_stage_inst_n28) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u21 ( .AN(ex_stage_inst_ex_alu_result[4]), 
        .B(rst), .Y(ex_stage_inst_n29) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u20 ( .AN(id_pipeline_reg_out[0]), .B(rst), 
        .Y(ex_stage_inst_n3) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u19 ( .AN(ex_stage_inst_ex_alu_result[5]), 
        .B(rst), .Y(ex_stage_inst_n30) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u18 ( .AN(ex_stage_inst_ex_alu_result[6]), 
        .B(rst), .Y(ex_stage_inst_n31) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u17 ( .AN(ex_stage_inst_ex_alu_result[7]), 
        .B(rst), .Y(ex_stage_inst_n32) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u16 ( .AN(ex_stage_inst_ex_alu_result[8]), 
        .B(rst), .Y(ex_stage_inst_n33) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u15 ( .AN(ex_stage_inst_ex_alu_result[9]), 
        .B(rst), .Y(ex_stage_inst_n34) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u14 ( .AN(ex_stage_inst_ex_alu_result[10]), 
        .B(rst), .Y(ex_stage_inst_n35) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u13 ( .AN(ex_stage_inst_ex_alu_result[11]), 
        .B(rst), .Y(ex_stage_inst_n36) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u12 ( .AN(ex_stage_inst_ex_alu_result[12]), 
        .B(rst), .Y(ex_stage_inst_n37) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u11 ( .AN(ex_stage_inst_ex_alu_result[13]), 
        .B(rst), .Y(ex_stage_inst_n38) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u10 ( .AN(ex_stage_inst_ex_alu_result[14]), 
        .B(rst), .Y(ex_stage_inst_n39) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u9 ( .AN(ex_op_dest[0]), .B(rst), .Y(
        ex_stage_inst_n4) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u8 ( .AN(ex_stage_inst_ex_alu_result[15]), 
        .B(rst), .Y(ex_stage_inst_n40) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u7 ( .AN(ex_op_dest[1]), .B(rst), .Y(
        ex_stage_inst_n5) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u6 ( .AN(ex_op_dest[2]), .B(rst), .Y(
        ex_stage_inst_n6) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u5 ( .AN(id_pipeline_reg_out[4]), .B(rst), 
        .Y(ex_stage_inst_n7) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u4 ( .AN(id_pipeline_reg_out[5]), .B(rst), 
        .Y(ex_stage_inst_n8) );
  NOR2B_X0P5M_A12TS ex_stage_inst_u3 ( .AN(id_pipeline_reg_out[6]), .B(rst), 
        .Y(ex_stage_inst_n9) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_24_ ( .D(ex_stage_inst_n27), .CK(clk), .Q(ex_pipeline_reg_out[24]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_25_ ( .D(ex_stage_inst_n28), .CK(clk), .Q(ex_pipeline_reg_out[25]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_5_ ( .D(ex_stage_inst_n8), 
        .CK(clk), .Q(ex_pipeline_reg_out[5]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_6_ ( .D(ex_stage_inst_n9), 
        .CK(clk), .Q(ex_pipeline_reg_out[6]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_7_ ( .D(ex_stage_inst_n10), 
        .CK(clk), .Q(ex_pipeline_reg_out[7]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_8_ ( .D(ex_stage_inst_n11), 
        .CK(clk), .Q(ex_pipeline_reg_out[8]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_9_ ( .D(ex_stage_inst_n12), 
        .CK(clk), .Q(ex_pipeline_reg_out[9]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_10_ ( .D(ex_stage_inst_n13), .CK(clk), .Q(ex_pipeline_reg_out[10]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_11_ ( .D(ex_stage_inst_n14), .CK(clk), .Q(ex_pipeline_reg_out[11]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_12_ ( .D(ex_stage_inst_n15), .CK(clk), .Q(ex_pipeline_reg_out[12]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_13_ ( .D(ex_stage_inst_n16), .CK(clk), .Q(ex_pipeline_reg_out[13]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_14_ ( .D(ex_stage_inst_n17), .CK(clk), .Q(ex_pipeline_reg_out[14]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_15_ ( .D(ex_stage_inst_n18), .CK(clk), .Q(ex_pipeline_reg_out[15]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_16_ ( .D(ex_stage_inst_n19), .CK(clk), .Q(ex_pipeline_reg_out[16]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_17_ ( .D(ex_stage_inst_n20), .CK(clk), .Q(ex_pipeline_reg_out[17]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_18_ ( .D(ex_stage_inst_n21), .CK(clk), .Q(ex_pipeline_reg_out[18]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_19_ ( .D(ex_stage_inst_n22), .CK(clk), .Q(ex_pipeline_reg_out[19]) );
  DFFQ_X3M_A12TS ex_stage_inst_pipeline_reg_out_reg_20_ ( .D(ex_stage_inst_n23), .CK(clk), .Q(ex_pipeline_reg_out[20]) );
  DFFQ_X2M_A12TS ex_stage_inst_pipeline_reg_out_reg_27_ ( .D(ex_stage_inst_n30), .CK(clk), .Q(ex_pipeline_reg_out[27]) );
  DFFQ_X2M_A12TS ex_stage_inst_pipeline_reg_out_reg_26_ ( .D(ex_stage_inst_n29), .CK(clk), .Q(ex_pipeline_reg_out[26]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_22_ ( .D(ex_stage_inst_n25), .CK(clk), .Q(ex_pipeline_reg_out[22]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_23_ ( .D(ex_stage_inst_n26), .CK(clk), .Q(ex_pipeline_reg_out[23]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_29_ ( .D(ex_stage_inst_n32), .CK(clk), .Q(ex_pipeline_reg_out[29]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_28_ ( .D(ex_stage_inst_n31), .CK(clk), .Q(ex_pipeline_reg_out[28]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_1_ ( .D(ex_stage_inst_n4), 
        .CK(clk), .Q(mem_op_dest[0]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_2_ ( .D(ex_stage_inst_n5), 
        .CK(clk), .Q(mem_op_dest[1]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_3_ ( .D(ex_stage_inst_n6), 
        .CK(clk), .Q(mem_op_dest[2]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_21_ ( .D(ex_stage_inst_n24), .CK(clk), .Q(ex_pipeline_reg_out[21]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_0_ ( .D(ex_stage_inst_n3), 
        .CK(clk), .Q(ex_pipeline_reg_out[0]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_4_ ( .D(ex_stage_inst_n7), 
        .CK(clk), .Q(ex_pipeline_reg_out[4]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_30_ ( .D(ex_stage_inst_n33), .CK(clk), .Q(ex_pipeline_reg_out[30]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_31_ ( .D(ex_stage_inst_n34), .CK(clk), .Q(ex_pipeline_reg_out[31]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_32_ ( .D(ex_stage_inst_n35), .CK(clk), .Q(ex_pipeline_reg_out[32]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_33_ ( .D(ex_stage_inst_n36), .CK(clk), .Q(ex_pipeline_reg_out[33]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_34_ ( .D(ex_stage_inst_n37), .CK(clk), .Q(ex_pipeline_reg_out[34]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_35_ ( .D(ex_stage_inst_n38), .CK(clk), .Q(ex_pipeline_reg_out[35]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_36_ ( .D(ex_stage_inst_n39), .CK(clk), .Q(ex_pipeline_reg_out[36]) );
  DFFQ_X1M_A12TS ex_stage_inst_pipeline_reg_out_reg_37_ ( .D(ex_stage_inst_n40), .CK(clk), .Q(ex_pipeline_reg_out[37]) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u226 ( .A(id_pipeline_reg_out[50]), 
        .Y(ex_stage_inst_alu_inst_n133) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u225 ( .A(id_pipeline_reg_out[22]), 
        .Y(ex_stage_inst_alu_inst_n209) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u224 ( .A(id_pipeline_reg_out[23]), 
        .Y(ex_stage_inst_alu_inst_n152) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u223 ( .A(
        ex_stage_inst_alu_inst_n209), .B(ex_stage_inst_alu_inst_n152), .Y(
        ex_stage_inst_alu_inst_n95) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u222 ( .A(ex_stage_inst_alu_inst_n95), 
        .Y(ex_stage_inst_alu_inst_n106) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u221 ( .A(id_pipeline_reg_out[53]), 
        .Y(ex_stage_inst_alu_inst_n34) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u220 ( .A(id_pipeline_reg_out[23]), 
        .B(id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_n96) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u219 ( .A(ex_stage_inst_alu_inst_n96), 
        .Y(ex_stage_inst_alu_inst_n107) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u218 ( .A(id_pipeline_reg_out[23]), 
        .B(ex_stage_inst_alu_inst_n209), .Y(ex_stage_inst_alu_inst_n116) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u217 ( .A(id_pipeline_reg_out[22]), 
        .B(ex_stage_inst_alu_inst_n152), .Y(ex_stage_inst_alu_inst_n117) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u216 ( .A0(
        ex_stage_inst_alu_inst_n116), .A1(id_pipeline_reg_out[52]), .B0(
        ex_stage_inst_alu_inst_n117), .B1(id_pipeline_reg_out[51]), .Y(
        ex_stage_inst_alu_inst_n208) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u215 ( .A0(
        ex_stage_inst_alu_inst_n133), .A1(ex_stage_inst_alu_inst_n106), .B0(
        ex_stage_inst_alu_inst_n34), .B1(ex_stage_inst_alu_inst_n107), .C0(
        ex_stage_inst_alu_inst_n208), .Y(ex_stage_inst_alu_inst_n31) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u214 ( .A(id_pipeline_reg_out[26]), 
        .Y(ex_stage_inst_alu_inst_n36) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u213 ( .A(id_pipeline_reg_out[25]), 
        .B(ex_stage_inst_alu_inst_n36), .Y(ex_stage_inst_alu_inst_n35) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u212 ( .A(ex_stage_inst_alu_inst_n35), 
        .Y(ex_stage_inst_alu_inst_n15) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u211 ( .A(
        ex_stage_inst_alu_inst_n15), .B(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_n73) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u210 ( .A(id_pipeline_reg_out[46]), 
        .Y(ex_stage_inst_alu_inst_n30) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u209 ( .A(id_pipeline_reg_out[49]), 
        .Y(ex_stage_inst_alu_inst_n188) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u208 ( .A0(
        ex_stage_inst_alu_inst_n116), .A1(id_pipeline_reg_out[48]), .B0(
        ex_stage_inst_alu_inst_n117), .B1(id_pipeline_reg_out[47]), .Y(
        ex_stage_inst_alu_inst_n207) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u207 ( .A0(
        ex_stage_inst_alu_inst_n30), .A1(ex_stage_inst_alu_inst_n106), .B0(
        ex_stage_inst_alu_inst_n188), .B1(ex_stage_inst_alu_inst_n107), .C0(
        ex_stage_inst_alu_inst_n207), .Y(ex_stage_inst_alu_inst_n32) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u206 ( .A(id_pipeline_reg_out[24]), 
        .Y(ex_stage_inst_alu_inst_n121) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u205 ( .A(
        ex_stage_inst_alu_inst_n15), .B(ex_stage_inst_alu_inst_n121), .Y(
        ex_stage_inst_alu_inst_n62) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u204 ( .A(id_pipeline_reg_out[26]), 
        .B(ex_stage_inst_alu_inst_n34), .Y(ex_stage_inst_alu_inst_n94) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u203 ( .A0(
        ex_stage_inst_alu_inst_n31), .A1(ex_stage_inst_alu_inst_n73), .B0(
        ex_stage_inst_alu_inst_n32), .B1(ex_stage_inst_alu_inst_n62), .C0(
        ex_stage_inst_alu_inst_n94), .Y(ex_stage_inst_alu_inst_n191) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u202 ( .A(id_pipeline_reg_out[38]), 
        .Y(ex_stage_inst_alu_inst_n200) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u201 ( .A(id_pipeline_reg_out[41]), 
        .Y(ex_stage_inst_alu_inst_n92) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u200 ( .A0(id_pipeline_reg_out[39]), 
        .A1(ex_stage_inst_alu_inst_n117), .B0(id_pipeline_reg_out[40]), .B1(
        ex_stage_inst_alu_inst_n116), .Y(ex_stage_inst_alu_inst_n206) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u199 ( .A0(
        ex_stage_inst_alu_inst_n106), .A1(ex_stage_inst_alu_inst_n200), .B0(
        ex_stage_inst_alu_inst_n107), .B1(ex_stage_inst_alu_inst_n92), .C0(
        ex_stage_inst_alu_inst_n206), .Y(ex_stage_inst_alu_inst_n201) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u198 ( .A(id_pipeline_reg_out[25]), 
        .Y(ex_stage_inst_alu_inst_n18) );
  NAND3_X0P5A_A12TS ex_stage_inst_alu_inst_u197 ( .A(
        ex_stage_inst_alu_inst_n18), .B(ex_stage_inst_alu_inst_n36), .C(
        ex_stage_inst_alu_inst_n121), .Y(ex_stage_inst_alu_inst_n42) );
  NAND3_X0P5A_A12TS ex_stage_inst_alu_inst_u196 ( .A(
        ex_stage_inst_alu_inst_n18), .B(ex_stage_inst_alu_inst_n36), .C(
        id_pipeline_reg_out[24]), .Y(ex_stage_inst_alu_inst_n49) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u195 ( .A(id_pipeline_reg_out[42]), 
        .Y(ex_stage_inst_alu_inst_n105) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u194 ( .A(id_pipeline_reg_out[45]), 
        .Y(ex_stage_inst_alu_inst_n51) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u193 ( .A(ex_stage_inst_alu_inst_n116), .Y(ex_stage_inst_alu_inst_n99) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u192 ( .A(ex_stage_inst_alu_inst_n117), .Y(ex_stage_inst_alu_inst_n100) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u191 ( .A0(id_pipeline_reg_out[44]), 
        .A1(ex_stage_inst_alu_inst_n99), .B0(id_pipeline_reg_out[43]), .B1(
        ex_stage_inst_alu_inst_n100), .Y(ex_stage_inst_alu_inst_n205) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u190 ( .A0(
        ex_stage_inst_alu_inst_n95), .A1(ex_stage_inst_alu_inst_n105), .B0(
        ex_stage_inst_alu_inst_n96), .B1(ex_stage_inst_alu_inst_n51), .C0(
        ex_stage_inst_alu_inst_n205), .Y(ex_stage_inst_alu_inst_n83) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u189 ( .A(id_pipeline_reg_out[56]), 
        .Y(ex_stage_inst_alu_inst_n196) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u188 ( .A(id_pipeline_reg_out[55]), 
        .Y(ex_stage_inst_alu_inst_n195) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u187 ( .A(id_pipeline_reg_out[32]), 
        .Y(ex_stage_inst_alu_inst_n189) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u186 ( .A(id_pipeline_reg_out[33]), 
        .Y(ex_stage_inst_alu_inst_n179) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u185 ( .A(id_pipeline_reg_out[34]), 
        .Y(ex_stage_inst_alu_inst_n168) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u184 ( .A(id_pipeline_reg_out[35]), 
        .Y(ex_stage_inst_alu_inst_n159) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u183 ( .A(
        ex_stage_inst_alu_inst_n189), .B(ex_stage_inst_alu_inst_n179), .C(
        ex_stage_inst_alu_inst_n168), .D(ex_stage_inst_alu_inst_n159), .Y(
        ex_stage_inst_alu_inst_n202) );
  OR4_X0P5M_A12TS ex_stage_inst_alu_inst_u182 ( .A(id_pipeline_reg_out[28]), 
        .B(id_pipeline_reg_out[29]), .C(id_pipeline_reg_out[30]), .D(
        id_pipeline_reg_out[31]), .Y(ex_stage_inst_alu_inst_n203) );
  OR3_X0P5M_A12TS ex_stage_inst_alu_inst_u181 ( .A(id_pipeline_reg_out[37]), 
        .B(id_pipeline_reg_out[27]), .C(id_pipeline_reg_out[36]), .Y(
        ex_stage_inst_alu_inst_n204) );
  OR6_X0P5M_A12TS ex_stage_inst_alu_inst_u180 ( .A(id_pipeline_reg_out[54]), 
        .B(ex_stage_inst_alu_inst_n196), .C(ex_stage_inst_alu_inst_n195), .D(
        ex_stage_inst_alu_inst_n202), .E(ex_stage_inst_alu_inst_n203), .F(
        ex_stage_inst_alu_inst_n204), .Y(ex_stage_inst_alu_inst_n2) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u179 ( .A(ex_stage_inst_alu_inst_n2), 
        .Y(ex_stage_inst_alu_inst_n44) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u178 ( .A0(
        ex_stage_inst_alu_inst_n201), .A1(ex_stage_inst_alu_inst_n42), .B0(
        ex_stage_inst_alu_inst_n49), .B1(ex_stage_inst_alu_inst_n83), .C0(
        ex_stage_inst_alu_inst_n44), .Y(ex_stage_inst_alu_inst_n192) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u177 ( .A(id_pipeline_reg_out[55]), 
        .B(ex_stage_inst_alu_inst_n196), .Y(ex_stage_inst_alu_inst_n14) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u176 ( .A(ex_stage_inst_alu_inst_n14), 
        .Y(ex_stage_inst_alu_inst_n149) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u175 ( .A(id_pipeline_reg_out[54]), 
        .B(ex_stage_inst_alu_inst_n149), .Y(ex_stage_inst_alu_inst_n12) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u174 ( .A(ex_stage_inst_alu_inst_n12), 
        .Y(ex_stage_inst_alu_inst_n8) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u173 ( .A(id_pipeline_reg_out[54]), 
        .Y(ex_stage_inst_alu_inst_n197) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u172 ( .A(
        ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(
        id_pipeline_reg_out[38]), .Y(ex_stage_inst_alu_inst_n198) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u171 ( .A0(
        id_pipeline_reg_out[22]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n200), .Y(
        ex_stage_inst_alu_inst_n199) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u170 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n198), .B0(
        id_pipeline_reg_out[22]), .C0(ex_stage_inst_alu_inst_n199), .Y(
        ex_stage_inst_alu_inst_n193) );
  NOR3_X0P5A_A12TS ex_stage_inst_alu_inst_u169 ( .A(
        ex_stage_inst_alu_inst_n196), .B(id_pipeline_reg_out[55]), .C(
        ex_stage_inst_alu_inst_n197), .Y(ex_stage_inst_alu_inst_n5) );
  NOR2_X0P5A_A12TS ex_stage_inst_alu_inst_u168 ( .A(id_pipeline_reg_out[55]), 
        .B(id_pipeline_reg_out[56]), .Y(ex_stage_inst_alu_inst_n6) );
  NOR3_X0P5A_A12TS ex_stage_inst_alu_inst_u167 ( .A(
        ex_stage_inst_alu_inst_n195), .B(ex_stage_inst_alu_inst_n196), .C(
        ex_stage_inst_alu_inst_n197), .Y(ex_stage_inst_alu_inst_n7) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u166 ( .A0(
        ex_stage_inst_alu_inst_n1130), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n490), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1450), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n194) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u165 ( .A0(
        ex_stage_inst_alu_inst_n191), .A1(ex_stage_inst_alu_inst_n192), .B0(
        ex_stage_inst_alu_inst_n193), .C0(ex_stage_inst_alu_inst_n194), .Y(
        ex_stage_inst_ex_alu_result[0]) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u164 ( .A(
        ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(
        id_pipeline_reg_out[48]), .Y(ex_stage_inst_alu_inst_n190) );
  OAI21_X0P5M_A12TS ex_stage_inst_alu_inst_u163 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n190), .B0(
        id_pipeline_reg_out[32]), .Y(ex_stage_inst_alu_inst_n181) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u162 ( .A(ex_stage_inst_alu_inst_n11), 
        .Y(ex_stage_inst_alu_inst_n84) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u161 ( .A0(
        ex_stage_inst_alu_inst_n84), .A1(ex_stage_inst_alu_inst_n189), .B0(
        ex_stage_inst_alu_inst_n8), .C0(id_pipeline_reg_out[48]), .Y(
        ex_stage_inst_alu_inst_n182) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u160 ( .A(id_pipeline_reg_out[52]), 
        .Y(ex_stage_inst_alu_inst_n163) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u159 ( .A(
        ex_stage_inst_alu_inst_n34), .B(ex_stage_inst_alu_inst_n163), .S0(
        ex_stage_inst_alu_inst_n106), .Y(ex_stage_inst_alu_inst_n61) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u158 ( .A(id_pipeline_reg_out[53]), 
        .B(ex_stage_inst_alu_inst_n18), .Y(ex_stage_inst_alu_inst_n37) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u157 ( .A(id_pipeline_reg_out[26]), 
        .B(ex_stage_inst_alu_inst_n37), .Y(ex_stage_inst_alu_inst_n75) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u156 ( .A(ex_stage_inst_alu_inst_n75), 
        .Y(ex_stage_inst_alu_inst_n47) );
  AOI31_X0P5M_A12TS ex_stage_inst_alu_inst_u155 ( .A0(id_pipeline_reg_out[24]), 
        .A1(id_pipeline_reg_out[23]), .A2(id_pipeline_reg_out[26]), .B0(
        ex_stage_inst_alu_inst_n47), .Y(ex_stage_inst_alu_inst_n185) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u154 ( .A(ex_stage_inst_alu_inst_n42), 
        .Y(ex_stage_inst_alu_inst_n21) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u153 ( .A0(
        ex_stage_inst_alu_inst_n99), .A1(ex_stage_inst_alu_inst_n133), .B0(
        ex_stage_inst_alu_inst_n100), .B1(ex_stage_inst_alu_inst_n188), .Y(
        ex_stage_inst_alu_inst_n187) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u152 ( .A0(id_pipeline_reg_out[48]), .A1(ex_stage_inst_alu_inst_n95), .B0(id_pipeline_reg_out[51]), .B1(
        ex_stage_inst_alu_inst_n96), .C0(ex_stage_inst_alu_inst_n187), .Y(
        ex_stage_inst_alu_inst_n122) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u151 ( .A0(
        ex_stage_inst_alu_inst_n21), .A1(ex_stage_inst_alu_inst_n122), .B0(
        id_pipeline_reg_out[25]), .B1(ex_stage_inst_alu_inst_n34), .C0(
        ex_stage_inst_alu_inst_n2), .Y(ex_stage_inst_alu_inst_n186) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u150 ( .A0(
        ex_stage_inst_alu_inst_n61), .A1(ex_stage_inst_alu_inst_n49), .B0(
        ex_stage_inst_alu_inst_n185), .C0(ex_stage_inst_alu_inst_n186), .Y(
        ex_stage_inst_alu_inst_n183) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u149 ( .A0(
        ex_stage_inst_alu_inst_n1230), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n590), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1550), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n184) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u148 ( .A(
        ex_stage_inst_alu_inst_n181), .B(ex_stage_inst_alu_inst_n182), .C(
        ex_stage_inst_alu_inst_n183), .D(ex_stage_inst_alu_inst_n184), .Y(
        ex_stage_inst_ex_alu_result[10]) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u147 ( .A(
        ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(
        id_pipeline_reg_out[49]), .Y(ex_stage_inst_alu_inst_n180) );
  OAI21_X0P5M_A12TS ex_stage_inst_alu_inst_u146 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n180), .B0(
        id_pipeline_reg_out[33]), .Y(ex_stage_inst_alu_inst_n172) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u145 ( .A0(
        ex_stage_inst_alu_inst_n84), .A1(ex_stage_inst_alu_inst_n179), .B0(
        ex_stage_inst_alu_inst_n8), .C0(id_pipeline_reg_out[49]), .Y(
        ex_stage_inst_alu_inst_n173) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u144 ( .A(id_pipeline_reg_out[51]), 
        .Y(ex_stage_inst_alu_inst_n162) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u143 ( .A0(
        ex_stage_inst_alu_inst_n162), .A1(ex_stage_inst_alu_inst_n116), .B0(
        ex_stage_inst_alu_inst_n133), .B1(ex_stage_inst_alu_inst_n117), .Y(
        ex_stage_inst_alu_inst_n178) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u142 ( .A0(
        ex_stage_inst_alu_inst_n106), .A1(id_pipeline_reg_out[49]), .B0(
        ex_stage_inst_alu_inst_n107), .B1(id_pipeline_reg_out[52]), .C0(
        ex_stage_inst_alu_inst_n178), .Y(ex_stage_inst_alu_inst_n46) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u141 ( .A(
        ex_stage_inst_alu_inst_n34), .B(ex_stage_inst_alu_inst_n46), .S0(
        ex_stage_inst_alu_inst_n21), .Y(ex_stage_inst_alu_inst_n176) );
  NOR2_X0P5A_A12TS ex_stage_inst_alu_inst_u140 ( .A(ex_stage_inst_alu_inst_n18), .B(ex_stage_inst_alu_inst_n36), .Y(ex_stage_inst_alu_inst_n81) );
  AOI31_X0P5M_A12TS ex_stage_inst_alu_inst_u139 ( .A0(id_pipeline_reg_out[24]), 
        .A1(ex_stage_inst_alu_inst_n95), .A2(id_pipeline_reg_out[26]), .B0(
        ex_stage_inst_alu_inst_n81), .Y(ex_stage_inst_alu_inst_n177) );
  NAND3_X0P5A_A12TS ex_stage_inst_alu_inst_u138 ( .A(
        ex_stage_inst_alu_inst_n176), .B(ex_stage_inst_alu_inst_n44), .C(
        ex_stage_inst_alu_inst_n177), .Y(ex_stage_inst_alu_inst_n174) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u137 ( .A0(
        ex_stage_inst_alu_inst_n1240), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n600), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1560), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n175) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u136 ( .A(
        ex_stage_inst_alu_inst_n172), .B(ex_stage_inst_alu_inst_n173), .C(
        ex_stage_inst_alu_inst_n174), .D(ex_stage_inst_alu_inst_n175), .Y(
        ex_stage_inst_ex_alu_result[11]) );
  NAND4B_X0P5M_A12TS ex_stage_inst_alu_inst_u135 ( .AN(
        ex_stage_inst_alu_inst_n37), .B(ex_stage_inst_alu_inst_n44), .C(
        id_pipeline_reg_out[26]), .D(ex_stage_inst_alu_inst_n121), .Y(
        ex_stage_inst_alu_inst_n153) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u134 ( .A0(
        id_pipeline_reg_out[26]), .A1(ex_stage_inst_alu_inst_n121), .B0(
        ex_stage_inst_alu_inst_n35), .C0(ex_stage_inst_alu_inst_n34), .Y(
        ex_stage_inst_alu_inst_n171) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u133 ( .A(
        ex_stage_inst_alu_inst_n171), .B(ex_stage_inst_alu_inst_n44), .Y(
        ex_stage_inst_alu_inst_n142) );
  NOR2_X0P5A_A12TS ex_stage_inst_alu_inst_u132 ( .A(ex_stage_inst_alu_inst_n2), 
        .B(ex_stage_inst_alu_inst_n42), .Y(ex_stage_inst_alu_inst_n150) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u131 ( .A0(
        id_pipeline_reg_out[34]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n133), .Y(
        ex_stage_inst_alu_inst_n170) );
  AOI21_X0P5M_A12TS ex_stage_inst_alu_inst_u130 ( .A0(
        ex_stage_inst_alu_inst_n150), .A1(ex_stage_inst_alu_inst_n31), .B0(
        ex_stage_inst_alu_inst_n170), .Y(ex_stage_inst_alu_inst_n164) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u129 ( .A(
        ex_stage_inst_alu_inst_n84), .B(ex_stage_inst_alu_inst_n149), .S0(
        id_pipeline_reg_out[50]), .Y(ex_stage_inst_alu_inst_n167) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u128 ( .A(
        ex_stage_inst_alu_inst_n610), .B(ex_stage_inst_alu_inst_n6), .Y(
        ex_stage_inst_alu_inst_n169) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u127 ( .A0(
        ex_stage_inst_alu_inst_n167), .A1(ex_stage_inst_alu_inst_n12), .B0(
        ex_stage_inst_alu_inst_n168), .C0(ex_stage_inst_alu_inst_n169), .Y(
        ex_stage_inst_alu_inst_n166) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u126 ( .A0(
        ex_stage_inst_alu_inst_n1570), .A1(ex_stage_inst_alu_inst_n7), .B0(
        ex_stage_inst_alu_inst_n1250), .B1(ex_stage_inst_alu_inst_n5), .C0(
        ex_stage_inst_alu_inst_n166), .Y(ex_stage_inst_alu_inst_n165) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u125 ( .A(
        ex_stage_inst_alu_inst_n153), .B(ex_stage_inst_alu_inst_n142), .C(
        ex_stage_inst_alu_inst_n164), .D(ex_stage_inst_alu_inst_n165), .Y(
        ex_stage_inst_ex_alu_result[12]) );
  NOR3_X0P5A_A12TS ex_stage_inst_alu_inst_u124 ( .A(
        ex_stage_inst_alu_inst_n107), .B(id_pipeline_reg_out[24]), .C(
        ex_stage_inst_alu_inst_n34), .Y(ex_stage_inst_alu_inst_n74) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u123 ( .A(
        ex_stage_inst_alu_inst_n74), .B(ex_stage_inst_alu_inst_n44), .C(
        id_pipeline_reg_out[26]), .D(ex_stage_inst_alu_inst_n18), .Y(
        ex_stage_inst_alu_inst_n154) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u122 ( .A0(
        ex_stage_inst_alu_inst_n162), .A1(ex_stage_inst_alu_inst_n106), .B0(
        ex_stage_inst_alu_inst_n163), .B1(ex_stage_inst_alu_inst_n100), .C0(
        ex_stage_inst_alu_inst_n34), .C1(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_n22) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u121 ( .A0(
        id_pipeline_reg_out[35]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n162), .Y(
        ex_stage_inst_alu_inst_n161) );
  AOI21_X0P5M_A12TS ex_stage_inst_alu_inst_u120 ( .A0(
        ex_stage_inst_alu_inst_n150), .A1(ex_stage_inst_alu_inst_n22), .B0(
        ex_stage_inst_alu_inst_n161), .Y(ex_stage_inst_alu_inst_n155) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u119 ( .A(
        ex_stage_inst_alu_inst_n84), .B(ex_stage_inst_alu_inst_n149), .S0(
        id_pipeline_reg_out[51]), .Y(ex_stage_inst_alu_inst_n158) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u118 ( .A(
        ex_stage_inst_alu_inst_n620), .B(ex_stage_inst_alu_inst_n6), .Y(
        ex_stage_inst_alu_inst_n160) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u117 ( .A0(
        ex_stage_inst_alu_inst_n158), .A1(ex_stage_inst_alu_inst_n12), .B0(
        ex_stage_inst_alu_inst_n159), .C0(ex_stage_inst_alu_inst_n160), .Y(
        ex_stage_inst_alu_inst_n157) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u116 ( .A0(
        ex_stage_inst_alu_inst_n1580), .A1(ex_stage_inst_alu_inst_n7), .B0(
        ex_stage_inst_alu_inst_n1260), .B1(ex_stage_inst_alu_inst_n5), .C0(
        ex_stage_inst_alu_inst_n157), .Y(ex_stage_inst_alu_inst_n156) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u115 ( .A(
        ex_stage_inst_alu_inst_n154), .B(ex_stage_inst_alu_inst_n142), .C(
        ex_stage_inst_alu_inst_n155), .D(ex_stage_inst_alu_inst_n156), .Y(
        ex_stage_inst_ex_alu_result[13]) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u114 ( .A(id_pipeline_reg_out[36]), 
        .Y(ex_stage_inst_alu_inst_n147) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u113 ( .A0(
        ex_stage_inst_alu_inst_n84), .A1(ex_stage_inst_alu_inst_n147), .B0(
        ex_stage_inst_alu_inst_n8), .C0(id_pipeline_reg_out[52]), .Y(
        ex_stage_inst_alu_inst_n141) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u112 ( .A(ex_stage_inst_alu_inst_n153), .Y(ex_stage_inst_alu_inst_n151) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u111 ( .A0(
        ex_stage_inst_alu_inst_n150), .A1(ex_stage_inst_alu_inst_n61), .B0(
        ex_stage_inst_alu_inst_n151), .B1(ex_stage_inst_alu_inst_n152), .Y(
        ex_stage_inst_alu_inst_n143) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u110 ( .A(
        ex_stage_inst_alu_inst_n84), .B(ex_stage_inst_alu_inst_n149), .S0(
        id_pipeline_reg_out[52]), .Y(ex_stage_inst_alu_inst_n146) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u109 ( .A(
        ex_stage_inst_alu_inst_n630), .B(ex_stage_inst_alu_inst_n6), .Y(
        ex_stage_inst_alu_inst_n148) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u108 ( .A0(
        ex_stage_inst_alu_inst_n146), .A1(ex_stage_inst_alu_inst_n12), .B0(
        ex_stage_inst_alu_inst_n147), .C0(ex_stage_inst_alu_inst_n148), .Y(
        ex_stage_inst_alu_inst_n145) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u107 ( .A0(
        ex_stage_inst_alu_inst_n1590), .A1(ex_stage_inst_alu_inst_n7), .B0(
        ex_stage_inst_alu_inst_n1270), .B1(ex_stage_inst_alu_inst_n5), .C0(
        ex_stage_inst_alu_inst_n145), .Y(ex_stage_inst_alu_inst_n144) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u106 ( .A(
        ex_stage_inst_alu_inst_n141), .B(ex_stage_inst_alu_inst_n142), .C(
        ex_stage_inst_alu_inst_n143), .D(ex_stage_inst_alu_inst_n144), .Y(
        ex_stage_inst_ex_alu_result[14]) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u105 ( .A(
        ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(
        id_pipeline_reg_out[37]), .Y(ex_stage_inst_alu_inst_n140) );
  AOI211_X0P5M_A12TS ex_stage_inst_alu_inst_u104 ( .A0(
        ex_stage_inst_alu_inst_n44), .A1(ex_stage_inst_alu_inst_n36), .B0(
        ex_stage_inst_alu_inst_n140), .C0(ex_stage_inst_alu_inst_n8), .Y(
        ex_stage_inst_alu_inst_n135) );
  NAND3_X0P5A_A12TS ex_stage_inst_alu_inst_u103 ( .A(id_pipeline_reg_out[53]), 
        .B(ex_stage_inst_alu_inst_n121), .C(ex_stage_inst_alu_inst_n106), .Y(
        ex_stage_inst_alu_inst_n48) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u102 ( .A(ex_stage_inst_alu_inst_n48), 
        .Y(ex_stage_inst_alu_inst_n138) );
  OAI21_X0P5M_A12TS ex_stage_inst_alu_inst_u101 ( .A0(id_pipeline_reg_out[53]), 
        .A1(ex_stage_inst_alu_inst_n11), .B0(ex_stage_inst_alu_inst_n12), .Y(
        ex_stage_inst_alu_inst_n139) );
  AOI32_X0P5M_A12TS ex_stage_inst_alu_inst_u100 ( .A0(
        ex_stage_inst_alu_inst_n44), .A1(ex_stage_inst_alu_inst_n18), .A2(
        ex_stage_inst_alu_inst_n138), .B0(id_pipeline_reg_out[37]), .B1(
        ex_stage_inst_alu_inst_n139), .Y(ex_stage_inst_alu_inst_n136) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u99 ( .A0(
        ex_stage_inst_alu_inst_n1280), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n640), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1600), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n137) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u98 ( .A0(
        ex_stage_inst_alu_inst_n135), .A1(ex_stage_inst_alu_inst_n34), .B0(
        ex_stage_inst_alu_inst_n136), .C0(ex_stage_inst_alu_inst_n137), .Y(
        ex_stage_inst_ex_alu_result[15]) );
  AOI21_X0P5M_A12TS ex_stage_inst_alu_inst_u97 ( .A0(
        ex_stage_inst_alu_inst_n107), .A1(id_pipeline_reg_out[24]), .B0(
        ex_stage_inst_alu_inst_n34), .Y(ex_stage_inst_alu_inst_n19) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u96 ( .A(id_pipeline_reg_out[47]), 
        .Y(ex_stage_inst_alu_inst_n13) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u95 ( .A0(
        ex_stage_inst_alu_inst_n116), .A1(id_pipeline_reg_out[49]), .B0(
        ex_stage_inst_alu_inst_n117), .B1(id_pipeline_reg_out[48]), .Y(
        ex_stage_inst_alu_inst_n134) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u94 ( .A0(
        ex_stage_inst_alu_inst_n13), .A1(ex_stage_inst_alu_inst_n106), .B0(
        ex_stage_inst_alu_inst_n133), .B1(ex_stage_inst_alu_inst_n107), .C0(
        ex_stage_inst_alu_inst_n134), .Y(ex_stage_inst_alu_inst_n20) );
  OAI222_X0P5M_A12TS ex_stage_inst_alu_inst_u93 ( .A0(
        ex_stage_inst_alu_inst_n22), .A1(ex_stage_inst_alu_inst_n73), .B0(
        ex_stage_inst_alu_inst_n19), .B1(ex_stage_inst_alu_inst_n75), .C0(
        ex_stage_inst_alu_inst_n20), .C1(ex_stage_inst_alu_inst_n62), .Y(
        ex_stage_inst_alu_inst_n123) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u92 ( .A(id_pipeline_reg_out[39]), 
        .Y(ex_stage_inst_alu_inst_n129) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u91 ( .A0(id_pipeline_reg_out[40]), 
        .A1(ex_stage_inst_alu_inst_n117), .B0(id_pipeline_reg_out[41]), .B1(
        ex_stage_inst_alu_inst_n116), .Y(ex_stage_inst_alu_inst_n132) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u90 ( .A0(
        ex_stage_inst_alu_inst_n106), .A1(ex_stage_inst_alu_inst_n129), .B0(
        ex_stage_inst_alu_inst_n107), .B1(ex_stage_inst_alu_inst_n105), .C0(
        ex_stage_inst_alu_inst_n132), .Y(ex_stage_inst_alu_inst_n130) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u89 ( .A(id_pipeline_reg_out[43]), 
        .Y(ex_stage_inst_alu_inst_n71) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u88 ( .A0(id_pipeline_reg_out[45]), 
        .A1(ex_stage_inst_alu_inst_n99), .B0(id_pipeline_reg_out[44]), .B1(
        ex_stage_inst_alu_inst_n100), .Y(ex_stage_inst_alu_inst_n131) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u87 ( .A0(
        ex_stage_inst_alu_inst_n95), .A1(ex_stage_inst_alu_inst_n71), .B0(
        ex_stage_inst_alu_inst_n96), .B1(ex_stage_inst_alu_inst_n30), .C0(
        ex_stage_inst_alu_inst_n131), .Y(ex_stage_inst_alu_inst_n72) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u86 ( .A0(
        ex_stage_inst_alu_inst_n130), .A1(ex_stage_inst_alu_inst_n42), .B0(
        ex_stage_inst_alu_inst_n49), .B1(ex_stage_inst_alu_inst_n72), .C0(
        ex_stage_inst_alu_inst_n44), .Y(ex_stage_inst_alu_inst_n124) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u85 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[39]), .Y(
        ex_stage_inst_alu_inst_n127) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u84 ( .A0(
        id_pipeline_reg_out[23]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n129), .Y(
        ex_stage_inst_alu_inst_n128) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u83 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n127), .B0(
        id_pipeline_reg_out[23]), .C0(ex_stage_inst_alu_inst_n128), .Y(
        ex_stage_inst_alu_inst_n125) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u82 ( .A0(
        ex_stage_inst_alu_inst_n1140), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n500), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1460), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n126) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u81 ( .A0(
        ex_stage_inst_alu_inst_n123), .A1(ex_stage_inst_alu_inst_n124), .B0(
        ex_stage_inst_alu_inst_n125), .C0(ex_stage_inst_alu_inst_n126), .Y(
        ex_stage_inst_ex_alu_result[1]) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u80 ( .A(ex_stage_inst_alu_inst_n122), 
        .Y(ex_stage_inst_alu_inst_n63) );
  NAND2_X0P5A_A12TS ex_stage_inst_alu_inst_u79 ( .A(ex_stage_inst_alu_inst_n81), .B(id_pipeline_reg_out[23]), .Y(ex_stage_inst_alu_inst_n64) );
  OA22_X0P5M_A12TS ex_stage_inst_alu_inst_u78 ( .A0(ex_stage_inst_alu_inst_n62), .A1(ex_stage_inst_alu_inst_n63), .B0(ex_stage_inst_alu_inst_n64), .B1(
        ex_stage_inst_alu_inst_n121), .Y(ex_stage_inst_alu_inst_n120) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u77 ( .A0(
        ex_stage_inst_alu_inst_n61), .A1(ex_stage_inst_alu_inst_n73), .B0(
        ex_stage_inst_alu_inst_n94), .C0(ex_stage_inst_alu_inst_n120), .Y(
        ex_stage_inst_alu_inst_n108) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u76 ( .A(id_pipeline_reg_out[40]), 
        .Y(ex_stage_inst_alu_inst_n114) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u75 ( .A0(id_pipeline_reg_out[41]), 
        .A1(ex_stage_inst_alu_inst_n117), .B0(id_pipeline_reg_out[42]), .B1(
        ex_stage_inst_alu_inst_n116), .Y(ex_stage_inst_alu_inst_n119) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u74 ( .A0(
        ex_stage_inst_alu_inst_n106), .A1(ex_stage_inst_alu_inst_n114), .B0(
        ex_stage_inst_alu_inst_n107), .B1(ex_stage_inst_alu_inst_n71), .C0(
        ex_stage_inst_alu_inst_n119), .Y(ex_stage_inst_alu_inst_n115) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u73 ( .A0(id_pipeline_reg_out[44]), 
        .A1(ex_stage_inst_alu_inst_n106), .B0(ex_stage_inst_alu_inst_n107), 
        .B1(id_pipeline_reg_out[47]), .Y(ex_stage_inst_alu_inst_n118) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u72 ( .A0(
        ex_stage_inst_alu_inst_n116), .A1(ex_stage_inst_alu_inst_n30), .B0(
        ex_stage_inst_alu_inst_n117), .B1(ex_stage_inst_alu_inst_n51), .C0(
        ex_stage_inst_alu_inst_n118), .Y(ex_stage_inst_alu_inst_n59) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u71 ( .A0(
        ex_stage_inst_alu_inst_n115), .A1(ex_stage_inst_alu_inst_n42), .B0(
        ex_stage_inst_alu_inst_n49), .B1(ex_stage_inst_alu_inst_n59), .C0(
        ex_stage_inst_alu_inst_n44), .Y(ex_stage_inst_alu_inst_n109) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u70 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[40]), .Y(
        ex_stage_inst_alu_inst_n112) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u69 ( .A0(
        id_pipeline_reg_out[24]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n114), .Y(
        ex_stage_inst_alu_inst_n113) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u68 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n112), .B0(
        id_pipeline_reg_out[24]), .C0(ex_stage_inst_alu_inst_n113), .Y(
        ex_stage_inst_alu_inst_n110) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u67 ( .A0(
        ex_stage_inst_alu_inst_n1150), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n510), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1470), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n111) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u66 ( .A0(
        ex_stage_inst_alu_inst_n108), .A1(ex_stage_inst_alu_inst_n109), .B0(
        ex_stage_inst_alu_inst_n110), .C0(ex_stage_inst_alu_inst_n111), .Y(
        ex_stage_inst_ex_alu_result[2]) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u65 ( .A(id_pipeline_reg_out[44]), 
        .Y(ex_stage_inst_alu_inst_n58) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u64 ( .A0(
        ex_stage_inst_alu_inst_n106), .A1(ex_stage_inst_alu_inst_n92), .B0(
        ex_stage_inst_alu_inst_n107), .B1(ex_stage_inst_alu_inst_n58), .Y(
        ex_stage_inst_alu_inst_n101) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u63 ( .A0(
        ex_stage_inst_alu_inst_n99), .A1(ex_stage_inst_alu_inst_n71), .B0(
        ex_stage_inst_alu_inst_n100), .B1(ex_stage_inst_alu_inst_n105), .Y(
        ex_stage_inst_alu_inst_n102) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u62 ( .A(ex_stage_inst_alu_inst_n62), 
        .Y(ex_stage_inst_alu_inst_n104) );
  AOI32_X0P5M_A12TS ex_stage_inst_alu_inst_u61 ( .A0(id_pipeline_reg_out[24]), 
        .A1(ex_stage_inst_alu_inst_n95), .A2(ex_stage_inst_alu_inst_n81), .B0(
        ex_stage_inst_alu_inst_n104), .B1(ex_stage_inst_alu_inst_n46), .Y(
        ex_stage_inst_alu_inst_n103) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u60 ( .A0(
        ex_stage_inst_alu_inst_n101), .A1(ex_stage_inst_alu_inst_n102), .B0(
        ex_stage_inst_alu_inst_n42), .C0(ex_stage_inst_alu_inst_n103), .Y(
        ex_stage_inst_alu_inst_n86) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u59 ( .A(id_pipeline_reg_out[48]), 
        .Y(ex_stage_inst_alu_inst_n97) );
  AOI22_X0P5M_A12TS ex_stage_inst_alu_inst_u58 ( .A0(
        ex_stage_inst_alu_inst_n99), .A1(id_pipeline_reg_out[47]), .B0(
        id_pipeline_reg_out[46]), .B1(ex_stage_inst_alu_inst_n100), .Y(
        ex_stage_inst_alu_inst_n98) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u57 ( .A0(
        ex_stage_inst_alu_inst_n95), .A1(ex_stage_inst_alu_inst_n51), .B0(
        ex_stage_inst_alu_inst_n96), .B1(ex_stage_inst_alu_inst_n97), .C0(
        ex_stage_inst_alu_inst_n98), .Y(ex_stage_inst_alu_inst_n43) );
  OAI21_X0P5M_A12TS ex_stage_inst_alu_inst_u56 ( .A0(id_pipeline_reg_out[53]), 
        .A1(ex_stage_inst_alu_inst_n73), .B0(ex_stage_inst_alu_inst_n94), .Y(
        ex_stage_inst_alu_inst_n82) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u55 ( .A(ex_stage_inst_alu_inst_n82), 
        .Y(ex_stage_inst_alu_inst_n93) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u54 ( .A0(
        ex_stage_inst_alu_inst_n49), .A1(ex_stage_inst_alu_inst_n43), .B0(
        ex_stage_inst_alu_inst_n44), .C0(ex_stage_inst_alu_inst_n93), .Y(
        ex_stage_inst_alu_inst_n87) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u53 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[41]), .Y(
        ex_stage_inst_alu_inst_n90) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u52 ( .A0(
        id_pipeline_reg_out[25]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n92), .Y(
        ex_stage_inst_alu_inst_n91) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u51 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n90), .B0(
        id_pipeline_reg_out[25]), .C0(ex_stage_inst_alu_inst_n91), .Y(
        ex_stage_inst_alu_inst_n88) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u50 ( .A0(
        ex_stage_inst_alu_inst_n1160), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n520), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1480), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n89) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u49 ( .A0(
        ex_stage_inst_alu_inst_n86), .A1(ex_stage_inst_alu_inst_n87), .B0(
        ex_stage_inst_alu_inst_n88), .C0(ex_stage_inst_alu_inst_n89), .Y(
        ex_stage_inst_ex_alu_result[3]) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u48 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[42]), .Y(
        ex_stage_inst_alu_inst_n85) );
  OAI21_X0P5M_A12TS ex_stage_inst_alu_inst_u47 ( .A0(ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n85), .B0(id_pipeline_reg_out[26]), .Y(
        ex_stage_inst_alu_inst_n76) );
  AO21A1AI2_X0P5M_A12TS ex_stage_inst_alu_inst_u46 ( .A0(
        ex_stage_inst_alu_inst_n84), .A1(ex_stage_inst_alu_inst_n36), .B0(
        ex_stage_inst_alu_inst_n8), .C0(id_pipeline_reg_out[42]), .Y(
        ex_stage_inst_alu_inst_n77) );
  OAI222_X0P5M_A12TS ex_stage_inst_alu_inst_u45 ( .A0(
        ex_stage_inst_alu_inst_n83), .A1(ex_stage_inst_alu_inst_n42), .B0(
        ex_stage_inst_alu_inst_n62), .B1(ex_stage_inst_alu_inst_n31), .C0(
        ex_stage_inst_alu_inst_n49), .C1(ex_stage_inst_alu_inst_n32), .Y(
        ex_stage_inst_alu_inst_n80) );
  AOI21_X0P5M_A12TS ex_stage_inst_alu_inst_u44 ( .A0(id_pipeline_reg_out[24]), 
        .A1(ex_stage_inst_alu_inst_n81), .B0(ex_stage_inst_alu_inst_n82), .Y(
        ex_stage_inst_alu_inst_n60) );
  NAND3B_X0P5M_A12TS ex_stage_inst_alu_inst_u43 ( .AN(
        ex_stage_inst_alu_inst_n80), .B(ex_stage_inst_alu_inst_n60), .C(
        ex_stage_inst_alu_inst_n44), .Y(ex_stage_inst_alu_inst_n78) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u42 ( .A0(
        ex_stage_inst_alu_inst_n1170), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n530), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1490), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n79) );
  NAND4_X0P5A_A12TS ex_stage_inst_alu_inst_u41 ( .A(ex_stage_inst_alu_inst_n76), .B(ex_stage_inst_alu_inst_n77), .C(ex_stage_inst_alu_inst_n78), .D(
        ex_stage_inst_alu_inst_n79), .Y(ex_stage_inst_ex_alu_result[4]) );
  OAI222_X0P5M_A12TS ex_stage_inst_alu_inst_u40 ( .A0(id_pipeline_reg_out[53]), 
        .A1(ex_stage_inst_alu_inst_n73), .B0(ex_stage_inst_alu_inst_n74), .B1(
        ex_stage_inst_alu_inst_n75), .C0(ex_stage_inst_alu_inst_n22), .C1(
        ex_stage_inst_alu_inst_n62), .Y(ex_stage_inst_alu_inst_n65) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u39 ( .A0(
        ex_stage_inst_alu_inst_n20), .A1(ex_stage_inst_alu_inst_n49), .B0(
        ex_stage_inst_alu_inst_n42), .B1(ex_stage_inst_alu_inst_n72), .C0(
        ex_stage_inst_alu_inst_n44), .Y(ex_stage_inst_alu_inst_n66) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u38 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[43]), .Y(
        ex_stage_inst_alu_inst_n69) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u37 ( .A0(
        id_pipeline_reg_out[27]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n71), .Y(
        ex_stage_inst_alu_inst_n70) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u36 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n69), .B0(
        id_pipeline_reg_out[27]), .C0(ex_stage_inst_alu_inst_n70), .Y(
        ex_stage_inst_alu_inst_n67) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u35 ( .A0(
        ex_stage_inst_alu_inst_n1180), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n540), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1500), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n68) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u34 ( .A0(
        ex_stage_inst_alu_inst_n65), .A1(ex_stage_inst_alu_inst_n66), .B0(
        ex_stage_inst_alu_inst_n67), .C0(ex_stage_inst_alu_inst_n68), .Y(
        ex_stage_inst_ex_alu_result[5]) );
  OAI221_X0P5M_A12TS ex_stage_inst_alu_inst_u33 ( .A0(
        ex_stage_inst_alu_inst_n61), .A1(ex_stage_inst_alu_inst_n62), .B0(
        ex_stage_inst_alu_inst_n63), .B1(ex_stage_inst_alu_inst_n49), .C0(
        ex_stage_inst_alu_inst_n64), .Y(ex_stage_inst_alu_inst_n52) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u32 ( .A0(
        ex_stage_inst_alu_inst_n42), .A1(ex_stage_inst_alu_inst_n59), .B0(
        ex_stage_inst_alu_inst_n44), .C0(ex_stage_inst_alu_inst_n60), .Y(
        ex_stage_inst_alu_inst_n53) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u31 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[44]), .Y(
        ex_stage_inst_alu_inst_n56) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u30 ( .A0(
        id_pipeline_reg_out[28]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n58), .Y(
        ex_stage_inst_alu_inst_n57) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u29 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n56), .B0(
        id_pipeline_reg_out[28]), .C0(ex_stage_inst_alu_inst_n57), .Y(
        ex_stage_inst_alu_inst_n54) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u28 ( .A0(
        ex_stage_inst_alu_inst_n1190), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n550), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1510), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n55) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u27 ( .A0(
        ex_stage_inst_alu_inst_n52), .A1(ex_stage_inst_alu_inst_n53), .B0(
        ex_stage_inst_alu_inst_n54), .C0(ex_stage_inst_alu_inst_n55), .Y(
        ex_stage_inst_ex_alu_result[6]) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u26 ( .A0(
        ex_stage_inst_alu_inst_n11), .A1(id_pipeline_reg_out[29]), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n51), .Y(
        ex_stage_inst_alu_inst_n38) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u25 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[45]), .Y(
        ex_stage_inst_alu_inst_n50) );
  OAI21_X0P5M_A12TS ex_stage_inst_alu_inst_u24 ( .A0(ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n50), .B0(id_pipeline_reg_out[29]), .Y(
        ex_stage_inst_alu_inst_n39) );
  INV_X0P5B_A12TS ex_stage_inst_alu_inst_u23 ( .A(ex_stage_inst_alu_inst_n49), 
        .Y(ex_stage_inst_alu_inst_n23) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u22 ( .A0(
        ex_stage_inst_alu_inst_n46), .A1(ex_stage_inst_alu_inst_n23), .B0(
        ex_stage_inst_alu_inst_n47), .B1(ex_stage_inst_alu_inst_n48), .C0(
        ex_stage_inst_alu_inst_n15), .C1(ex_stage_inst_alu_inst_n34), .Y(
        ex_stage_inst_alu_inst_n45) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u21 ( .A0(
        ex_stage_inst_alu_inst_n42), .A1(ex_stage_inst_alu_inst_n43), .B0(
        ex_stage_inst_alu_inst_n44), .C0(ex_stage_inst_alu_inst_n45), .Y(
        ex_stage_inst_alu_inst_n40) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u20 ( .A0(
        ex_stage_inst_alu_inst_n1200), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n560), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1520), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n41) );
  NAND4B_X0P5M_A12TS ex_stage_inst_alu_inst_u19 ( .AN(
        ex_stage_inst_alu_inst_n38), .B(ex_stage_inst_alu_inst_n39), .C(
        ex_stage_inst_alu_inst_n40), .D(ex_stage_inst_alu_inst_n41), .Y(
        ex_stage_inst_ex_alu_result[7]) );
  OAI22_X0P5M_A12TS ex_stage_inst_alu_inst_u18 ( .A0(
        ex_stage_inst_alu_inst_n34), .A1(ex_stage_inst_alu_inst_n35), .B0(
        ex_stage_inst_alu_inst_n36), .B1(ex_stage_inst_alu_inst_n37), .Y(
        ex_stage_inst_alu_inst_n33) );
  AOI221_X0P5M_A12TS ex_stage_inst_alu_inst_u17 ( .A0(
        ex_stage_inst_alu_inst_n31), .A1(ex_stage_inst_alu_inst_n23), .B0(
        ex_stage_inst_alu_inst_n32), .B1(ex_stage_inst_alu_inst_n21), .C0(
        ex_stage_inst_alu_inst_n33), .Y(ex_stage_inst_alu_inst_n24) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u16 ( .A(ex_stage_inst_alu_inst_n11), .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[46]), .Y(
        ex_stage_inst_alu_inst_n28) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u15 ( .A0(
        id_pipeline_reg_out[30]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n30), .Y(
        ex_stage_inst_alu_inst_n29) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u14 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n28), .B0(
        id_pipeline_reg_out[30]), .C0(ex_stage_inst_alu_inst_n29), .Y(
        ex_stage_inst_alu_inst_n25) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u13 ( .A0(
        ex_stage_inst_alu_inst_n1210), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n570), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1530), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n27) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u12 ( .A0(
        ex_stage_inst_alu_inst_n24), .A1(ex_stage_inst_alu_inst_n2), .B0(
        ex_stage_inst_alu_inst_n25), .C0(ex_stage_inst_alu_inst_n27), .Y(
        ex_stage_inst_ex_alu_result[8]) );
  AO22_X0P5M_A12TS ex_stage_inst_alu_inst_u11 ( .A0(ex_stage_inst_alu_inst_n20), .A1(ex_stage_inst_alu_inst_n21), .B0(ex_stage_inst_alu_inst_n22), .B1(
        ex_stage_inst_alu_inst_n23), .Y(ex_stage_inst_alu_inst_n16) );
  AND3_X0P5M_A12TS ex_stage_inst_alu_inst_u10 ( .A(id_pipeline_reg_out[26]), 
        .B(ex_stage_inst_alu_inst_n18), .C(ex_stage_inst_alu_inst_n19), .Y(
        ex_stage_inst_alu_inst_n17) );
  AOI211_X0P5M_A12TS ex_stage_inst_alu_inst_u9 ( .A0(
        ex_stage_inst_alu_inst_n15), .A1(id_pipeline_reg_out[53]), .B0(
        ex_stage_inst_alu_inst_n16), .C0(ex_stage_inst_alu_inst_n17), .Y(
        ex_stage_inst_alu_inst_n1) );
  MXIT2_X0P5M_A12TS ex_stage_inst_alu_inst_u8 ( .A(ex_stage_inst_alu_inst_n11), 
        .B(ex_stage_inst_alu_inst_n14), .S0(id_pipeline_reg_out[47]), .Y(
        ex_stage_inst_alu_inst_n9) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u7 ( .A0(
        id_pipeline_reg_out[31]), .A1(ex_stage_inst_alu_inst_n11), .B0(
        ex_stage_inst_alu_inst_n12), .C0(ex_stage_inst_alu_inst_n13), .Y(
        ex_stage_inst_alu_inst_n10) );
  OA21A1OI2_X0P5M_A12TS ex_stage_inst_alu_inst_u6 ( .A0(
        ex_stage_inst_alu_inst_n8), .A1(ex_stage_inst_alu_inst_n9), .B0(
        id_pipeline_reg_out[31]), .C0(ex_stage_inst_alu_inst_n10), .Y(
        ex_stage_inst_alu_inst_n3) );
  AOI222_X0P5M_A12TS ex_stage_inst_alu_inst_u5 ( .A0(
        ex_stage_inst_alu_inst_n1220), .A1(ex_stage_inst_alu_inst_n5), .B0(
        ex_stage_inst_alu_inst_n580), .B1(ex_stage_inst_alu_inst_n6), .C0(
        ex_stage_inst_alu_inst_n1540), .C1(ex_stage_inst_alu_inst_n7), .Y(
        ex_stage_inst_alu_inst_n4) );
  OAI211_X0P5M_A12TS ex_stage_inst_alu_inst_u4 ( .A0(ex_stage_inst_alu_inst_n1), .A1(ex_stage_inst_alu_inst_n2), .B0(ex_stage_inst_alu_inst_n3), .C0(
        ex_stage_inst_alu_inst_n4), .Y(ex_stage_inst_ex_alu_result[9]) );
  TIELO_X1M_A12TS ex_stage_inst_alu_inst_u3 ( .Y(ex_stage_inst_alu_inst_n26)
         );
  NAND3_X1M_A12TS ex_stage_inst_alu_inst_u2 ( .A(ex_stage_inst_alu_inst_n197), 
        .B(ex_stage_inst_alu_inst_n195), .C(id_pipeline_reg_out[56]), .Y(
        ex_stage_inst_alu_inst_n11) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u16 ( .A(
        id_pipeline_reg_out[22]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[0]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u15 ( .A(
        id_pipeline_reg_out[32]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[10]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u14 ( .A(
        id_pipeline_reg_out[33]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[11]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u13 ( .A(
        id_pipeline_reg_out[34]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[12]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u12 ( .A(
        id_pipeline_reg_out[35]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[13]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u11 ( .A(
        id_pipeline_reg_out[36]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[14]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u10 ( .A(
        id_pipeline_reg_out[37]), .B(id_pipeline_reg_out[54]), .Y(
        ex_stage_inst_alu_inst_r316_b_as[15]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u9 ( .A(id_pipeline_reg_out[23]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[1]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u8 ( .A(id_pipeline_reg_out[24]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[2]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u7 ( .A(id_pipeline_reg_out[25]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[3]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u6 ( .A(id_pipeline_reg_out[26]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[4]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u5 ( .A(id_pipeline_reg_out[27]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[5]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u4 ( .A(id_pipeline_reg_out[28]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[6]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u3 ( .A(id_pipeline_reg_out[29]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[7]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u2 ( .A(id_pipeline_reg_out[30]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[8]) );
  XOR2_X0P5M_A12TS ex_stage_inst_alu_inst_r316_u1 ( .A(id_pipeline_reg_out[31]), .B(id_pipeline_reg_out[54]), .Y(ex_stage_inst_alu_inst_r316_b_as[9]) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_0 ( .A(id_pipeline_reg_out[38]), .B(ex_stage_inst_alu_inst_r316_b_as[0]), .CI(id_pipeline_reg_out[54]), .CO(
        ex_stage_inst_alu_inst_r316_carry_1_), .S(ex_stage_inst_alu_inst_n490)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_1 ( .A(id_pipeline_reg_out[39]), .B(ex_stage_inst_alu_inst_r316_b_as[1]), .CI(
        ex_stage_inst_alu_inst_r316_carry_1_), .CO(
        ex_stage_inst_alu_inst_r316_carry_2_), .S(ex_stage_inst_alu_inst_n500)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_2 ( .A(id_pipeline_reg_out[40]), .B(ex_stage_inst_alu_inst_r316_b_as[2]), .CI(
        ex_stage_inst_alu_inst_r316_carry_2_), .CO(
        ex_stage_inst_alu_inst_r316_carry_3_), .S(ex_stage_inst_alu_inst_n510)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_3 ( .A(id_pipeline_reg_out[41]), .B(ex_stage_inst_alu_inst_r316_b_as[3]), .CI(
        ex_stage_inst_alu_inst_r316_carry_3_), .CO(
        ex_stage_inst_alu_inst_r316_carry_4_), .S(ex_stage_inst_alu_inst_n520)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_4 ( .A(id_pipeline_reg_out[42]), .B(ex_stage_inst_alu_inst_r316_b_as[4]), .CI(
        ex_stage_inst_alu_inst_r316_carry_4_), .CO(
        ex_stage_inst_alu_inst_r316_carry_5_), .S(ex_stage_inst_alu_inst_n530)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_5 ( .A(id_pipeline_reg_out[43]), .B(ex_stage_inst_alu_inst_r316_b_as[5]), .CI(
        ex_stage_inst_alu_inst_r316_carry_5_), .CO(
        ex_stage_inst_alu_inst_r316_carry_6_), .S(ex_stage_inst_alu_inst_n540)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_6 ( .A(id_pipeline_reg_out[44]), .B(ex_stage_inst_alu_inst_r316_b_as[6]), .CI(
        ex_stage_inst_alu_inst_r316_carry_6_), .CO(
        ex_stage_inst_alu_inst_r316_carry_7_), .S(ex_stage_inst_alu_inst_n550)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_7 ( .A(id_pipeline_reg_out[45]), .B(ex_stage_inst_alu_inst_r316_b_as[7]), .CI(
        ex_stage_inst_alu_inst_r316_carry_7_), .CO(
        ex_stage_inst_alu_inst_r316_carry_8_), .S(ex_stage_inst_alu_inst_n560)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_8 ( .A(id_pipeline_reg_out[46]), .B(ex_stage_inst_alu_inst_r316_b_as[8]), .CI(
        ex_stage_inst_alu_inst_r316_carry_8_), .CO(
        ex_stage_inst_alu_inst_r316_carry_9_), .S(ex_stage_inst_alu_inst_n570)
         );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_9 ( .A(id_pipeline_reg_out[47]), .B(ex_stage_inst_alu_inst_r316_b_as[9]), .CI(
        ex_stage_inst_alu_inst_r316_carry_9_), .CO(
        ex_stage_inst_alu_inst_r316_carry_10_), .S(ex_stage_inst_alu_inst_n580) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_10 ( .A(
        id_pipeline_reg_out[48]), .B(ex_stage_inst_alu_inst_r316_b_as[10]), 
        .CI(ex_stage_inst_alu_inst_r316_carry_10_), .CO(
        ex_stage_inst_alu_inst_r316_carry_11_), .S(ex_stage_inst_alu_inst_n590) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_11 ( .A(
        id_pipeline_reg_out[49]), .B(ex_stage_inst_alu_inst_r316_b_as[11]), 
        .CI(ex_stage_inst_alu_inst_r316_carry_11_), .CO(
        ex_stage_inst_alu_inst_r316_carry_12_), .S(ex_stage_inst_alu_inst_n600) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_12 ( .A(
        id_pipeline_reg_out[50]), .B(ex_stage_inst_alu_inst_r316_b_as[12]), 
        .CI(ex_stage_inst_alu_inst_r316_carry_12_), .CO(
        ex_stage_inst_alu_inst_r316_carry_13_), .S(ex_stage_inst_alu_inst_n610) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_13 ( .A(
        id_pipeline_reg_out[51]), .B(ex_stage_inst_alu_inst_r316_b_as[13]), 
        .CI(ex_stage_inst_alu_inst_r316_carry_13_), .CO(
        ex_stage_inst_alu_inst_r316_carry_14_), .S(ex_stage_inst_alu_inst_n620) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_14 ( .A(
        id_pipeline_reg_out[52]), .B(ex_stage_inst_alu_inst_r316_b_as[14]), 
        .CI(ex_stage_inst_alu_inst_r316_carry_14_), .CO(
        ex_stage_inst_alu_inst_r316_carry_15_), .S(ex_stage_inst_alu_inst_n630) );
  ADDF_X1M_A12TS ex_stage_inst_alu_inst_r316_u1_15 ( .A(
        id_pipeline_reg_out[53]), .B(ex_stage_inst_alu_inst_r316_b_as[15]), 
        .CI(ex_stage_inst_alu_inst_r316_carry_15_), .CO(), .S(
        ex_stage_inst_alu_inst_n640) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u216 ( .A(
        id_pipeline_reg_out[31]), .B(id_pipeline_reg_out[32]), .Y(
        ex_stage_inst_alu_inst_sll_36_n146) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u215 ( .A(
        id_pipeline_reg_out[35]), .B(id_pipeline_reg_out[36]), .Y(
        ex_stage_inst_alu_inst_sll_36_n145) );
  NAND2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u214 ( .A(
        ex_stage_inst_alu_inst_sll_36_n145), .B(
        ex_stage_inst_alu_inst_sll_36_n146), .Y(
        ex_stage_inst_alu_inst_sll_36_n86) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u213 ( .A(
        id_pipeline_reg_out[29]), .B(id_pipeline_reg_out[30]), .Y(
        ex_stage_inst_alu_inst_sll_36_n89) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u212 ( .A(
        ex_stage_inst_alu_inst_sll_36_n89), .B(id_pipeline_reg_out[37]), .Y(
        ex_stage_inst_alu_inst_sll_36_n87) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u211 ( .A(
        id_pipeline_reg_out[28]), .B(id_pipeline_reg_out[27]), .Y(
        ex_stage_inst_alu_inst_sll_36_n88) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u210 ( .A(
        ex_stage_inst_alu_inst_sll_36_n63), .B(
        ex_stage_inst_alu_inst_sll_36_n59), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n47) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u209 ( .A(
        ex_stage_inst_alu_inst_sll_36_n47), .B(
        ex_stage_inst_alu_inst_sll_36_n39), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n31) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u208 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n31), .Y(
        ex_stage_inst_alu_inst_sll_36_n15) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u207 ( .A(
        ex_stage_inst_alu_inst_sll_36_n15), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1250) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u206 ( .A(
        ex_stage_inst_alu_inst_sll_36_n82), .B(
        ex_stage_inst_alu_inst_sll_36_n80), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n66) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u205 ( .A(
        ex_stage_inst_alu_inst_sll_36_n66), .B(
        ex_stage_inst_alu_inst_sll_36_n62), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n50) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u204 ( .A(
        ex_stage_inst_alu_inst_sll_36_n50), .B(
        ex_stage_inst_alu_inst_sll_36_n42), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n34) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u203 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n34), .Y(
        ex_stage_inst_alu_inst_sll_36_n18) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u202 ( .A(
        ex_stage_inst_alu_inst_sll_36_n81), .B(
        ex_stage_inst_alu_inst_sll_36_n79), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n65) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u201 ( .A(
        ex_stage_inst_alu_inst_sll_36_n65), .B(
        ex_stage_inst_alu_inst_sll_36_n61), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n49) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u200 ( .A(
        ex_stage_inst_alu_inst_sll_36_n49), .B(
        ex_stage_inst_alu_inst_sll_36_n41), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n33) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u199 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n33), .Y(
        ex_stage_inst_alu_inst_sll_36_n17) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u198 ( .A(
        ex_stage_inst_alu_inst_sll_36_n80), .B(
        ex_stage_inst_alu_inst_sll_36_n78), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n64) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u197 ( .A(
        ex_stage_inst_alu_inst_sll_36_n64), .B(
        ex_stage_inst_alu_inst_sll_36_n60), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n48) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u196 ( .A(
        ex_stage_inst_alu_inst_sll_36_n48), .B(
        ex_stage_inst_alu_inst_sll_36_n40), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n32) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u195 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n32), .Y(
        ex_stage_inst_alu_inst_sll_36_n16) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u194 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_sll_36_n52), .Y(
        ex_stage_inst_alu_inst_sll_36_n36) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u193 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_sll_36_n51), .Y(
        ex_stage_inst_alu_inst_sll_36_n35) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u192 ( .BN(
        id_pipeline_reg_out[22]), .A(id_pipeline_reg_out[38]), .Y(
        ex_stage_inst_alu_inst_sll_36_n67) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u191 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_sll_36_n54), .Y(
        ex_stage_inst_alu_inst_sll_36_n38) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u190 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_sll_36_n53), .Y(
        ex_stage_inst_alu_inst_sll_36_n37) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u189 ( .A(
        id_pipeline_reg_out[53]), .B(id_pipeline_reg_out[52]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n82) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u188 ( .A(
        id_pipeline_reg_out[52]), .B(id_pipeline_reg_out[51]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n81) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u187 ( .A(
        ex_stage_inst_alu_inst_sll_36_n79), .B(
        ex_stage_inst_alu_inst_sll_36_n77), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n63) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u186 ( .A(
        ex_stage_inst_alu_inst_sll_36_n68), .B(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n52) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u185 ( .A(
        ex_stage_inst_alu_inst_sll_36_n67), .B(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n51) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u184 ( .A(
        id_pipeline_reg_out[33]), .B(id_pipeline_reg_out[34]), .Y(
        ex_stage_inst_alu_inst_sll_36_n91) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u183 ( .A(
        ex_stage_inst_alu_inst_sll_36_n86), .B(
        ex_stage_inst_alu_inst_sll_36_n87), .Y(
        ex_stage_inst_alu_inst_sll_36_n84) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u182 ( .A(
        ex_stage_inst_alu_inst_sll_36_n88), .B(
        ex_stage_inst_alu_inst_sll_36_n91), .Y(
        ex_stage_inst_alu_inst_sll_36_n85) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u181 ( .A(
        ex_stage_inst_alu_inst_sll_36_n42), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n26) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u180 ( .A(
        ex_stage_inst_alu_inst_sll_36_n41), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n25) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u179 ( .A(
        ex_stage_inst_alu_inst_sll_36_n40), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n24) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u178 ( .A(
        ex_stage_inst_alu_inst_sll_36_n39), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n23) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u177 ( .A(
        ex_stage_inst_alu_inst_sll_36_n38), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n22) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u176 ( .A(
        ex_stage_inst_alu_inst_sll_36_n37), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n21) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u175 ( .A(
        ex_stage_inst_alu_inst_sll_36_n36), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n20) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u174 ( .A(
        ex_stage_inst_alu_inst_sll_36_n35), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n19) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u173 ( .A(
        id_pipeline_reg_out[51]), .B(id_pipeline_reg_out[50]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n80) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u172 ( .A(
        id_pipeline_reg_out[49]), .B(id_pipeline_reg_out[48]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n78) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u171 ( .A(
        id_pipeline_reg_out[47]), .B(id_pipeline_reg_out[46]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n76) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u170 ( .A(
        id_pipeline_reg_out[45]), .B(id_pipeline_reg_out[44]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n74) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u169 ( .A(
        id_pipeline_reg_out[43]), .B(id_pipeline_reg_out[42]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n72) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u168 ( .A(
        id_pipeline_reg_out[41]), .B(id_pipeline_reg_out[40]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n70) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u167 ( .A(
        id_pipeline_reg_out[50]), .B(id_pipeline_reg_out[49]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n79) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u166 ( .A(
        id_pipeline_reg_out[48]), .B(id_pipeline_reg_out[47]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n77) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u165 ( .A(
        id_pipeline_reg_out[46]), .B(id_pipeline_reg_out[45]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n75) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u164 ( .A(
        id_pipeline_reg_out[44]), .B(id_pipeline_reg_out[43]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n73) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u163 ( .A(
        id_pipeline_reg_out[42]), .B(id_pipeline_reg_out[41]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n71) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u162 ( .A(
        id_pipeline_reg_out[40]), .B(id_pipeline_reg_out[39]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n69) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u161 ( .A(
        ex_stage_inst_alu_inst_sll_36_n78), .B(
        ex_stage_inst_alu_inst_sll_36_n76), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n62) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u160 ( .A(
        ex_stage_inst_alu_inst_sll_36_n74), .B(
        ex_stage_inst_alu_inst_sll_36_n72), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n58) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u159 ( .A(
        ex_stage_inst_alu_inst_sll_36_n77), .B(
        ex_stage_inst_alu_inst_sll_36_n75), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n61) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u158 ( .A(
        ex_stage_inst_alu_inst_sll_36_n73), .B(
        ex_stage_inst_alu_inst_sll_36_n71), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n57) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u157 ( .A(
        ex_stage_inst_alu_inst_sll_36_n76), .B(
        ex_stage_inst_alu_inst_sll_36_n74), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n60) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u156 ( .A(
        ex_stage_inst_alu_inst_sll_36_n72), .B(
        ex_stage_inst_alu_inst_sll_36_n70), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n56) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u155 ( .A(
        ex_stage_inst_alu_inst_sll_36_n75), .B(
        ex_stage_inst_alu_inst_sll_36_n73), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n59) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u154 ( .A(
        ex_stage_inst_alu_inst_sll_36_n71), .B(
        ex_stage_inst_alu_inst_sll_36_n69), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n55) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u153 ( .A(
        ex_stage_inst_alu_inst_sll_36_n58), .B(
        ex_stage_inst_alu_inst_sll_36_n54), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n42) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u152 ( .A(
        ex_stage_inst_alu_inst_sll_36_n57), .B(
        ex_stage_inst_alu_inst_sll_36_n53), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n41) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u151 ( .A(
        ex_stage_inst_alu_inst_sll_36_n56), .B(
        ex_stage_inst_alu_inst_sll_36_n52), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n40) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u150 ( .A(
        ex_stage_inst_alu_inst_sll_36_n55), .B(
        ex_stage_inst_alu_inst_sll_36_n51), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n39) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u149 ( .A(
        id_pipeline_reg_out[39]), .B(id_pipeline_reg_out[38]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_sll_36_n68) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u148 ( .A(
        ex_stage_inst_alu_inst_sll_36_n62), .B(
        ex_stage_inst_alu_inst_sll_36_n58), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n46) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u147 ( .A(
        ex_stage_inst_alu_inst_sll_36_n46), .B(
        ex_stage_inst_alu_inst_sll_36_n38), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n30) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u146 ( .A(
        ex_stage_inst_alu_inst_sll_36_n61), .B(
        ex_stage_inst_alu_inst_sll_36_n57), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n45) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u145 ( .A(
        ex_stage_inst_alu_inst_sll_36_n45), .B(
        ex_stage_inst_alu_inst_sll_36_n37), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n29) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u144 ( .A(
        ex_stage_inst_alu_inst_sll_36_n60), .B(
        ex_stage_inst_alu_inst_sll_36_n56), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n44) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u143 ( .A(
        ex_stage_inst_alu_inst_sll_36_n44), .B(
        ex_stage_inst_alu_inst_sll_36_n36), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n28) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u142 ( .A(
        ex_stage_inst_alu_inst_sll_36_n59), .B(
        ex_stage_inst_alu_inst_sll_36_n55), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_sll_36_n43) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u141 ( .A(
        ex_stage_inst_alu_inst_sll_36_n43), .B(
        ex_stage_inst_alu_inst_sll_36_n35), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_sll_36_n27) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u140 ( .A(
        ex_stage_inst_alu_inst_sll_36_n70), .B(
        ex_stage_inst_alu_inst_sll_36_n68), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n54) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_sll_36_u139 ( .A(
        ex_stage_inst_alu_inst_sll_36_n69), .B(
        ex_stage_inst_alu_inst_sll_36_n67), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_sll_36_n53) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u138 ( .A(
        ex_stage_inst_alu_inst_sll_36_n18), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1280) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u137 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n28), .Y(
        ex_stage_inst_alu_inst_sll_36_n12) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u136 ( .A(
        ex_stage_inst_alu_inst_sll_36_n12), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1220) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u135 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n27), .Y(
        ex_stage_inst_alu_inst_sll_36_n11) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u134 ( .A(
        ex_stage_inst_alu_inst_sll_36_n11), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1210) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u133 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n25), .Y(
        ex_stage_inst_alu_inst_sll_36_n9) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u132 ( .A(
        ex_stage_inst_alu_inst_sll_36_n9), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1190) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u131 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n24), .Y(
        ex_stage_inst_alu_inst_sll_36_n8) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u130 ( .A(
        ex_stage_inst_alu_inst_sll_36_n8), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1180) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u129 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n22), .Y(
        ex_stage_inst_alu_inst_sll_36_n6) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u128 ( .A(
        ex_stage_inst_alu_inst_sll_36_n6), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1160) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u127 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n21), .Y(
        ex_stage_inst_alu_inst_sll_36_n5) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u126 ( .A(
        ex_stage_inst_alu_inst_sll_36_n5), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1150) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u125 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n20), .Y(
        ex_stage_inst_alu_inst_sll_36_n4) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u124 ( .A(
        ex_stage_inst_alu_inst_sll_36_n4), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1140) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u123 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n19), .Y(
        ex_stage_inst_alu_inst_sll_36_n3) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u122 ( .A(
        ex_stage_inst_alu_inst_sll_36_n3), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1130) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u121 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n30), .Y(
        ex_stage_inst_alu_inst_sll_36_n14) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u120 ( .A(
        ex_stage_inst_alu_inst_sll_36_n14), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1240) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u119 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n29), .Y(
        ex_stage_inst_alu_inst_sll_36_n13) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u118 ( .A(
        ex_stage_inst_alu_inst_sll_36_n13), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1230) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u117 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n23), .Y(
        ex_stage_inst_alu_inst_sll_36_n7) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u116 ( .A(
        ex_stage_inst_alu_inst_sll_36_n7), .B(ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1170) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u115 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_sll_36_n26), .Y(
        ex_stage_inst_alu_inst_sll_36_n10) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u114 ( .A(
        ex_stage_inst_alu_inst_sll_36_n10), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1200) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u113 ( .A(
        ex_stage_inst_alu_inst_sll_36_n17), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1270) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_sll_36_u112 ( .A(
        ex_stage_inst_alu_inst_sll_36_n16), .B(
        ex_stage_inst_alu_inst_sll_36_n2), .Y(ex_stage_inst_alu_inst_n1260) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_sll_36_u111 ( .A(
        ex_stage_inst_alu_inst_sll_36_n84), .B(
        ex_stage_inst_alu_inst_sll_36_n85), .Y(
        ex_stage_inst_alu_inst_sll_36_n2) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u217 ( .A(
        id_pipeline_reg_out[31]), .B(id_pipeline_reg_out[32]), .Y(
        ex_stage_inst_alu_inst_srl_40_n148) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u216 ( .A(
        id_pipeline_reg_out[35]), .B(id_pipeline_reg_out[36]), .Y(
        ex_stage_inst_alu_inst_srl_40_n147) );
  NAND2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u215 ( .A(
        ex_stage_inst_alu_inst_srl_40_n147), .B(
        ex_stage_inst_alu_inst_srl_40_n148), .Y(
        ex_stage_inst_alu_inst_srl_40_n86) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u214 ( .A(
        id_pipeline_reg_out[29]), .B(id_pipeline_reg_out[30]), .Y(
        ex_stage_inst_alu_inst_srl_40_n89) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u213 ( .A(
        ex_stage_inst_alu_inst_srl_40_n89), .B(id_pipeline_reg_out[37]), .Y(
        ex_stage_inst_alu_inst_srl_40_n87) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u212 ( .A(
        id_pipeline_reg_out[28]), .B(id_pipeline_reg_out[27]), .Y(
        ex_stage_inst_alu_inst_srl_40_n88) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u211 ( .A(
        ex_stage_inst_alu_inst_srl_40_n47), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n31) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u210 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n31), .Y(
        ex_stage_inst_alu_inst_srl_40_n15) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u209 ( .A(
        ex_stage_inst_alu_inst_srl_40_n15), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1570) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u208 ( .A(
        ex_stage_inst_alu_inst_srl_40_n50), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n34) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u207 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n34), .Y(
        ex_stage_inst_alu_inst_srl_40_n18) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u206 ( .A(
        ex_stage_inst_alu_inst_srl_40_n49), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n33) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u205 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n33), .Y(
        ex_stage_inst_alu_inst_srl_40_n17) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u204 ( .A(
        ex_stage_inst_alu_inst_srl_40_n48), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n32) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u203 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n32), .Y(
        ex_stage_inst_alu_inst_srl_40_n16) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u202 ( .A(
        ex_stage_inst_alu_inst_srl_40_n46), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n30) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u201 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n30), .Y(
        ex_stage_inst_alu_inst_srl_40_n14) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u200 ( .A(
        ex_stage_inst_alu_inst_srl_40_n45), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n29) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u199 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n29), .Y(
        ex_stage_inst_alu_inst_srl_40_n13) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u198 ( .A(
        ex_stage_inst_alu_inst_srl_40_n44), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n28) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u197 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n28), .Y(
        ex_stage_inst_alu_inst_srl_40_n12) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u196 ( .A(
        ex_stage_inst_alu_inst_srl_40_n43), .B(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n27) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u195 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n27), .Y(
        ex_stage_inst_alu_inst_srl_40_n11) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u194 ( .A(
        ex_stage_inst_alu_inst_srl_40_n58), .B(
        ex_stage_inst_alu_inst_srl_40_n62), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n42) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u193 ( .A(
        ex_stage_inst_alu_inst_srl_40_n42), .B(
        ex_stage_inst_alu_inst_srl_40_n50), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n26) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u192 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n26), .Y(
        ex_stage_inst_alu_inst_srl_40_n10) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u191 ( .A(
        ex_stage_inst_alu_inst_srl_40_n57), .B(
        ex_stage_inst_alu_inst_srl_40_n61), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n41) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u190 ( .A(
        ex_stage_inst_alu_inst_srl_40_n41), .B(
        ex_stage_inst_alu_inst_srl_40_n49), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n25) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u189 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n25), .Y(
        ex_stage_inst_alu_inst_srl_40_n9) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u188 ( .A(
        ex_stage_inst_alu_inst_srl_40_n56), .B(
        ex_stage_inst_alu_inst_srl_40_n60), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n40) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u187 ( .A(
        ex_stage_inst_alu_inst_srl_40_n40), .B(
        ex_stage_inst_alu_inst_srl_40_n48), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n24) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u186 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n24), .Y(
        ex_stage_inst_alu_inst_srl_40_n8) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u185 ( .A(
        ex_stage_inst_alu_inst_srl_40_n55), .B(
        ex_stage_inst_alu_inst_srl_40_n59), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n39) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u184 ( .A(
        ex_stage_inst_alu_inst_srl_40_n39), .B(
        ex_stage_inst_alu_inst_srl_40_n47), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n23) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u183 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n23), .Y(
        ex_stage_inst_alu_inst_srl_40_n7) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u182 ( .A(
        ex_stage_inst_alu_inst_srl_40_n70), .B(
        ex_stage_inst_alu_inst_srl_40_n72), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n54) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u181 ( .A(
        ex_stage_inst_alu_inst_srl_40_n54), .B(
        ex_stage_inst_alu_inst_srl_40_n58), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n38) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u180 ( .A(
        ex_stage_inst_alu_inst_srl_40_n38), .B(
        ex_stage_inst_alu_inst_srl_40_n46), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n22) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u179 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n22), .Y(
        ex_stage_inst_alu_inst_srl_40_n6) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u178 ( .A(
        ex_stage_inst_alu_inst_srl_40_n69), .B(
        ex_stage_inst_alu_inst_srl_40_n71), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n53) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u177 ( .A(
        ex_stage_inst_alu_inst_srl_40_n53), .B(
        ex_stage_inst_alu_inst_srl_40_n57), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n37) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u176 ( .A(
        ex_stage_inst_alu_inst_srl_40_n37), .B(
        ex_stage_inst_alu_inst_srl_40_n45), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n21) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u175 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n21), .Y(
        ex_stage_inst_alu_inst_srl_40_n5) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u174 ( .A(
        ex_stage_inst_alu_inst_srl_40_n68), .B(
        ex_stage_inst_alu_inst_srl_40_n70), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n52) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u173 ( .A(
        ex_stage_inst_alu_inst_srl_40_n52), .B(
        ex_stage_inst_alu_inst_srl_40_n56), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n36) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u172 ( .A(
        ex_stage_inst_alu_inst_srl_40_n36), .B(
        ex_stage_inst_alu_inst_srl_40_n44), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n20) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u171 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n20), .Y(
        ex_stage_inst_alu_inst_srl_40_n4) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u170 ( .A(
        ex_stage_inst_alu_inst_srl_40_n67), .B(
        ex_stage_inst_alu_inst_srl_40_n69), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n51) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u169 ( .A(
        ex_stage_inst_alu_inst_srl_40_n51), .B(
        ex_stage_inst_alu_inst_srl_40_n55), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n35) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u168 ( .A(
        ex_stage_inst_alu_inst_srl_40_n35), .B(
        ex_stage_inst_alu_inst_srl_40_n43), .S0(id_pipeline_reg_out[25]), .Y(
        ex_stage_inst_alu_inst_srl_40_n19) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u167 ( .BN(
        id_pipeline_reg_out[26]), .A(ex_stage_inst_alu_inst_srl_40_n19), .Y(
        ex_stage_inst_alu_inst_srl_40_n3) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u166 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_srl_40_n66), .Y(
        ex_stage_inst_alu_inst_srl_40_n50) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u165 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_srl_40_n65), .Y(
        ex_stage_inst_alu_inst_srl_40_n49) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u164 ( .BN(
        id_pipeline_reg_out[22]), .A(id_pipeline_reg_out[53]), .Y(
        ex_stage_inst_alu_inst_srl_40_n82) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u163 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_srl_40_n64), .Y(
        ex_stage_inst_alu_inst_srl_40_n48) );
  NAND2XB_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u162 ( .BN(
        id_pipeline_reg_out[24]), .A(ex_stage_inst_alu_inst_srl_40_n63), .Y(
        ex_stage_inst_alu_inst_srl_40_n47) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u161 ( .A(
        id_pipeline_reg_out[39]), .B(id_pipeline_reg_out[40]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n68) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u160 ( .A(
        id_pipeline_reg_out[38]), .B(id_pipeline_reg_out[39]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n67) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u159 ( .A(
        ex_stage_inst_alu_inst_srl_40_n82), .B(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n66) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u158 ( .A(
        ex_stage_inst_alu_inst_srl_40_n81), .B(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n65) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u157 ( .A(
        id_pipeline_reg_out[33]), .B(id_pipeline_reg_out[34]), .Y(
        ex_stage_inst_alu_inst_srl_40_n91) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u156 ( .A(
        ex_stage_inst_alu_inst_srl_40_n86), .B(
        ex_stage_inst_alu_inst_srl_40_n87), .Y(
        ex_stage_inst_alu_inst_srl_40_n84) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u155 ( .A(
        ex_stage_inst_alu_inst_srl_40_n88), .B(
        ex_stage_inst_alu_inst_srl_40_n91), .Y(
        ex_stage_inst_alu_inst_srl_40_n85) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u154 ( .A(
        id_pipeline_reg_out[51]), .B(id_pipeline_reg_out[52]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n80) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u153 ( .A(
        id_pipeline_reg_out[50]), .B(id_pipeline_reg_out[51]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n79) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u152 ( .A(
        id_pipeline_reg_out[49]), .B(id_pipeline_reg_out[50]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n78) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u151 ( .A(
        id_pipeline_reg_out[48]), .B(id_pipeline_reg_out[49]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n77) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u150 ( .A(
        id_pipeline_reg_out[47]), .B(id_pipeline_reg_out[48]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n76) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u149 ( .A(
        id_pipeline_reg_out[46]), .B(id_pipeline_reg_out[47]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n75) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u148 ( .A(
        id_pipeline_reg_out[45]), .B(id_pipeline_reg_out[46]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n74) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u147 ( .A(
        id_pipeline_reg_out[44]), .B(id_pipeline_reg_out[45]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n73) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u146 ( .A(
        id_pipeline_reg_out[43]), .B(id_pipeline_reg_out[44]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n72) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u145 ( .A(
        id_pipeline_reg_out[42]), .B(id_pipeline_reg_out[43]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n71) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u144 ( .A(
        id_pipeline_reg_out[41]), .B(id_pipeline_reg_out[42]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n70) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u143 ( .A(
        id_pipeline_reg_out[40]), .B(id_pipeline_reg_out[41]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n69) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u142 ( .A(
        ex_stage_inst_alu_inst_srl_40_n78), .B(
        ex_stage_inst_alu_inst_srl_40_n80), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n62) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u141 ( .A(
        ex_stage_inst_alu_inst_srl_40_n77), .B(
        ex_stage_inst_alu_inst_srl_40_n79), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n61) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u140 ( .A(
        ex_stage_inst_alu_inst_srl_40_n76), .B(
        ex_stage_inst_alu_inst_srl_40_n78), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n60) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u139 ( .A(
        ex_stage_inst_alu_inst_srl_40_n75), .B(
        ex_stage_inst_alu_inst_srl_40_n77), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n59) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u138 ( .A(
        ex_stage_inst_alu_inst_srl_40_n74), .B(
        ex_stage_inst_alu_inst_srl_40_n76), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n58) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u137 ( .A(
        ex_stage_inst_alu_inst_srl_40_n73), .B(
        ex_stage_inst_alu_inst_srl_40_n75), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n57) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u136 ( .A(
        ex_stage_inst_alu_inst_srl_40_n72), .B(
        ex_stage_inst_alu_inst_srl_40_n74), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n56) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u135 ( .A(
        ex_stage_inst_alu_inst_srl_40_n71), .B(
        ex_stage_inst_alu_inst_srl_40_n73), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n55) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u134 ( .A(
        ex_stage_inst_alu_inst_srl_40_n62), .B(
        ex_stage_inst_alu_inst_srl_40_n66), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n46) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u133 ( .A(
        ex_stage_inst_alu_inst_srl_40_n61), .B(
        ex_stage_inst_alu_inst_srl_40_n65), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n45) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u132 ( .A(
        ex_stage_inst_alu_inst_srl_40_n60), .B(
        ex_stage_inst_alu_inst_srl_40_n64), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n44) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u131 ( .A(
        ex_stage_inst_alu_inst_srl_40_n59), .B(
        ex_stage_inst_alu_inst_srl_40_n63), .S0(id_pipeline_reg_out[24]), .Y(
        ex_stage_inst_alu_inst_srl_40_n43) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u130 ( .A(
        id_pipeline_reg_out[52]), .B(id_pipeline_reg_out[53]), .S0(
        id_pipeline_reg_out[22]), .Y(ex_stage_inst_alu_inst_srl_40_n81) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u129 ( .A(
        ex_stage_inst_alu_inst_srl_40_n80), .B(
        ex_stage_inst_alu_inst_srl_40_n82), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n64) );
  MXIT2_X0P7M_A12TS ex_stage_inst_alu_inst_srl_40_u128 ( .A(
        ex_stage_inst_alu_inst_srl_40_n79), .B(
        ex_stage_inst_alu_inst_srl_40_n81), .S0(id_pipeline_reg_out[23]), .Y(
        ex_stage_inst_alu_inst_srl_40_n63) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u127 ( .A(
        ex_stage_inst_alu_inst_srl_40_n18), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1600) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u126 ( .A(
        ex_stage_inst_alu_inst_srl_40_n12), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1540) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u125 ( .A(
        ex_stage_inst_alu_inst_srl_40_n11), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1530) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u124 ( .A(
        ex_stage_inst_alu_inst_srl_40_n9), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1510) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u123 ( .A(
        ex_stage_inst_alu_inst_srl_40_n8), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1500) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u122 ( .A(
        ex_stage_inst_alu_inst_srl_40_n6), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1480) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u121 ( .A(
        ex_stage_inst_alu_inst_srl_40_n5), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1470) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u120 ( .A(
        ex_stage_inst_alu_inst_srl_40_n4), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1460) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u119 ( .A(
        ex_stage_inst_alu_inst_srl_40_n3), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1450) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u118 ( .A(
        ex_stage_inst_alu_inst_srl_40_n14), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1560) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u117 ( .A(
        ex_stage_inst_alu_inst_srl_40_n13), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1550) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u116 ( .A(
        ex_stage_inst_alu_inst_srl_40_n7), .B(ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1490) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u115 ( .A(
        ex_stage_inst_alu_inst_srl_40_n10), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1520) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u114 ( .A(
        ex_stage_inst_alu_inst_srl_40_n17), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1590) );
  NOR2_X1A_A12TS ex_stage_inst_alu_inst_srl_40_u113 ( .A(
        ex_stage_inst_alu_inst_srl_40_n16), .B(
        ex_stage_inst_alu_inst_srl_40_n2), .Y(ex_stage_inst_alu_inst_n1580) );
  OR2_X1M_A12TS ex_stage_inst_alu_inst_srl_40_u112 ( .A(
        ex_stage_inst_alu_inst_srl_40_n84), .B(
        ex_stage_inst_alu_inst_srl_40_n85), .Y(
        ex_stage_inst_alu_inst_srl_40_n2) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u39 ( .AN(mem_stage_inst_mem_read_data[2]), 
        .B(rst), .Y(mem_stage_inst_n10) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u38 ( .AN(mem_stage_inst_mem_read_data[3]), 
        .B(rst), .Y(mem_stage_inst_n11) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u37 ( .AN(mem_stage_inst_mem_read_data[4]), 
        .B(rst), .Y(mem_stage_inst_n12) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u36 ( .AN(mem_stage_inst_mem_read_data[5]), 
        .B(rst), .Y(mem_stage_inst_n13) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u35 ( .AN(mem_stage_inst_mem_read_data[6]), 
        .B(rst), .Y(mem_stage_inst_n14) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u34 ( .AN(mem_stage_inst_mem_read_data[7]), 
        .B(rst), .Y(mem_stage_inst_n15) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u33 ( .AN(mem_stage_inst_mem_read_data[8]), 
        .B(rst), .Y(mem_stage_inst_n16) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u32 ( .AN(mem_stage_inst_mem_read_data[9]), 
        .B(rst), .Y(mem_stage_inst_n17) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u31 ( .AN(mem_stage_inst_mem_read_data[10]), 
        .B(rst), .Y(mem_stage_inst_n18) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u30 ( .AN(mem_stage_inst_mem_read_data[11]), 
        .B(rst), .Y(mem_stage_inst_n19) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u29 ( .AN(mem_stage_inst_mem_read_data[12]), 
        .B(rst), .Y(mem_stage_inst_n20) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u28 ( .AN(mem_stage_inst_mem_read_data[13]), 
        .B(rst), .Y(mem_stage_inst_n21) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u27 ( .AN(mem_stage_inst_mem_read_data[14]), 
        .B(rst), .Y(mem_stage_inst_n22) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u26 ( .AN(mem_stage_inst_mem_read_data[15]), 
        .B(rst), .Y(mem_stage_inst_n23) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u25 ( .AN(ex_pipeline_reg_out[22]), .B(rst), 
        .Y(mem_stage_inst_n24) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u24 ( .AN(ex_pipeline_reg_out[23]), .B(rst), 
        .Y(mem_stage_inst_n25) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u23 ( .AN(ex_pipeline_reg_out[24]), .B(rst), 
        .Y(mem_stage_inst_n26) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u22 ( .AN(ex_pipeline_reg_out[25]), .B(rst), 
        .Y(mem_stage_inst_n27) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u21 ( .AN(ex_pipeline_reg_out[26]), .B(rst), 
        .Y(mem_stage_inst_n28) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u20 ( .AN(ex_pipeline_reg_out[27]), .B(rst), 
        .Y(mem_stage_inst_n29) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u19 ( .AN(ex_pipeline_reg_out[0]), .B(rst), 
        .Y(mem_stage_inst_n3) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u18 ( .AN(ex_pipeline_reg_out[28]), .B(rst), 
        .Y(mem_stage_inst_n30) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u17 ( .AN(ex_pipeline_reg_out[29]), .B(rst), 
        .Y(mem_stage_inst_n31) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u16 ( .AN(ex_pipeline_reg_out[30]), .B(rst), 
        .Y(mem_stage_inst_n32) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u15 ( .AN(ex_pipeline_reg_out[31]), .B(rst), 
        .Y(mem_stage_inst_n33) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u14 ( .AN(ex_pipeline_reg_out[32]), .B(rst), 
        .Y(mem_stage_inst_n34) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u13 ( .AN(ex_pipeline_reg_out[33]), .B(rst), 
        .Y(mem_stage_inst_n35) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u12 ( .AN(ex_pipeline_reg_out[34]), .B(rst), 
        .Y(mem_stage_inst_n36) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u11 ( .AN(ex_pipeline_reg_out[35]), .B(rst), 
        .Y(mem_stage_inst_n37) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u10 ( .AN(ex_pipeline_reg_out[36]), .B(rst), 
        .Y(mem_stage_inst_n38) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u9 ( .AN(ex_pipeline_reg_out[37]), .B(rst), 
        .Y(mem_stage_inst_n39) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u8 ( .AN(mem_op_dest[0]), .B(rst), .Y(
        mem_stage_inst_n4) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u7 ( .AN(mem_op_dest[1]), .B(rst), .Y(
        mem_stage_inst_n5) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u6 ( .AN(mem_op_dest[2]), .B(rst), .Y(
        mem_stage_inst_n6) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u5 ( .AN(ex_pipeline_reg_out[4]), .B(rst), 
        .Y(mem_stage_inst_n7) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u4 ( .AN(mem_stage_inst_mem_read_data[0]), 
        .B(rst), .Y(mem_stage_inst_n8) );
  NOR2B_X0P5M_A12TS mem_stage_inst_u3 ( .AN(mem_stage_inst_mem_read_data[1]), 
        .B(rst), .Y(mem_stage_inst_n9) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_0_ ( .D(mem_stage_inst_n3), .CK(clk), .Q(mem_pipeline_reg_out[0]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_2_ ( .D(mem_stage_inst_n5), .CK(clk), .Q(reg_write_dest[1]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_1_ ( .D(mem_stage_inst_n4), .CK(clk), .Q(reg_write_dest[0]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_3_ ( .D(mem_stage_inst_n6), .CK(clk), .Q(reg_write_dest[2]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_4_ ( .D(mem_stage_inst_n7), .CK(clk), .Q(reg_write_en) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_5_ ( .D(mem_stage_inst_n8), .CK(clk), .Q(mem_pipeline_reg_out[5]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_6_ ( .D(mem_stage_inst_n9), .CK(clk), .Q(mem_pipeline_reg_out[6]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_7_ ( .D(
        mem_stage_inst_n10), .CK(clk), .Q(mem_pipeline_reg_out[7]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_8_ ( .D(
        mem_stage_inst_n11), .CK(clk), .Q(mem_pipeline_reg_out[8]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_9_ ( .D(
        mem_stage_inst_n12), .CK(clk), .Q(mem_pipeline_reg_out[9]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_10_ ( .D(
        mem_stage_inst_n13), .CK(clk), .Q(mem_pipeline_reg_out[10]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_11_ ( .D(
        mem_stage_inst_n14), .CK(clk), .Q(mem_pipeline_reg_out[11]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_12_ ( .D(
        mem_stage_inst_n15), .CK(clk), .Q(mem_pipeline_reg_out[12]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_13_ ( .D(
        mem_stage_inst_n16), .CK(clk), .Q(mem_pipeline_reg_out[13]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_14_ ( .D(
        mem_stage_inst_n17), .CK(clk), .Q(mem_pipeline_reg_out[14]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_15_ ( .D(
        mem_stage_inst_n18), .CK(clk), .Q(mem_pipeline_reg_out[15]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_16_ ( .D(
        mem_stage_inst_n19), .CK(clk), .Q(mem_pipeline_reg_out[16]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_17_ ( .D(
        mem_stage_inst_n20), .CK(clk), .Q(mem_pipeline_reg_out[17]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_18_ ( .D(
        mem_stage_inst_n21), .CK(clk), .Q(mem_pipeline_reg_out[18]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_19_ ( .D(
        mem_stage_inst_n22), .CK(clk), .Q(mem_pipeline_reg_out[19]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_20_ ( .D(
        mem_stage_inst_n23), .CK(clk), .Q(mem_pipeline_reg_out[20]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_21_ ( .D(
        mem_stage_inst_n24), .CK(clk), .Q(mem_pipeline_reg_out[21]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_22_ ( .D(
        mem_stage_inst_n25), .CK(clk), .Q(mem_pipeline_reg_out[22]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_23_ ( .D(
        mem_stage_inst_n26), .CK(clk), .Q(mem_pipeline_reg_out[23]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_24_ ( .D(
        mem_stage_inst_n27), .CK(clk), .Q(mem_pipeline_reg_out[24]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_25_ ( .D(
        mem_stage_inst_n28), .CK(clk), .Q(mem_pipeline_reg_out[25]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_26_ ( .D(
        mem_stage_inst_n29), .CK(clk), .Q(mem_pipeline_reg_out[26]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_27_ ( .D(
        mem_stage_inst_n30), .CK(clk), .Q(mem_pipeline_reg_out[27]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_28_ ( .D(
        mem_stage_inst_n31), .CK(clk), .Q(mem_pipeline_reg_out[28]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_29_ ( .D(
        mem_stage_inst_n32), .CK(clk), .Q(mem_pipeline_reg_out[29]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_30_ ( .D(
        mem_stage_inst_n33), .CK(clk), .Q(mem_pipeline_reg_out[30]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_31_ ( .D(
        mem_stage_inst_n34), .CK(clk), .Q(mem_pipeline_reg_out[31]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_32_ ( .D(
        mem_stage_inst_n35), .CK(clk), .Q(mem_pipeline_reg_out[32]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_33_ ( .D(
        mem_stage_inst_n36), .CK(clk), .Q(mem_pipeline_reg_out[33]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_34_ ( .D(
        mem_stage_inst_n37), .CK(clk), .Q(mem_pipeline_reg_out[34]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_35_ ( .D(
        mem_stage_inst_n38), .CK(clk), .Q(mem_pipeline_reg_out[35]) );
  DFFQ_X1M_A12TS mem_stage_inst_pipeline_reg_out_reg_36_ ( .D(
        mem_stage_inst_n39), .CK(clk), .Q(mem_pipeline_reg_out[36]) );
  NOR2B_X0P5M_A12TS mem_stage_inst_dmem_u5986 ( .AN(ex_pipeline_reg_out[21]), 
        .B(ex_pipeline_reg_out[29]), .Y(mem_stage_inst_dmem_n5926) );
  INV_X0P5B_A12TS mem_stage_inst_dmem_u5985 ( .A(ex_pipeline_reg_out[28]), .Y(
        mem_stage_inst_dmem_n5856) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5984 ( .A(mem_stage_inst_dmem_n5926), 
        .B(mem_stage_inst_dmem_n5856), .Y(mem_stage_inst_dmem_n5713) );
  INV_X0P5B_A12TS mem_stage_inst_dmem_u5983 ( .A(ex_pipeline_reg_out[26]), .Y(
        mem_stage_inst_dmem_n5965) );
  NOR2_X0P5A_A12TS mem_stage_inst_dmem_u5982 ( .A(mem_stage_inst_dmem_n5965), 
        .B(ex_pipeline_reg_out[27]), .Y(mem_stage_inst_dmem_n5768) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5981 ( .A(mem_stage_inst_dmem_n5713), 
        .B(mem_stage_inst_dmem_n5768), .Y(mem_stage_inst_dmem_n5669) );
  NOR2_X0P5A_A12TS mem_stage_inst_dmem_u5980 ( .A(mem_stage_inst_dmem_n218), 
        .B(mem_stage_inst_dmem_n66), .Y(mem_stage_inst_dmem_n5953) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5979 ( .A(mem_stage_inst_dmem_n5953), 
        .B(mem_stage_inst_dmem_n204), .C(mem_stage_inst_dmem_n164), .Y(
        mem_stage_inst_dmem_n5700) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5978 ( .A(mem_stage_inst_dmem_n5669), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5666) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5977 ( .A(
        mem_stage_inst_dmem_ram_27__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1000) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5976 ( .A(
        mem_stage_inst_dmem_ram_27__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1001) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5975 ( .A(
        mem_stage_inst_dmem_ram_27__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1002) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5974 ( .A(
        mem_stage_inst_dmem_ram_27__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1003) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5973 ( .A(
        mem_stage_inst_dmem_ram_27__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1004) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5972 ( .A(
        mem_stage_inst_dmem_ram_27__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1005) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5971 ( .A(
        mem_stage_inst_dmem_ram_27__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1006) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5970 ( .A(
        mem_stage_inst_dmem_ram_27__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1007) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5969 ( .A(
        mem_stage_inst_dmem_ram_27__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1008) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5968 ( .A(
        mem_stage_inst_dmem_ram_27__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1009) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5967 ( .A(
        mem_stage_inst_dmem_ram_27__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1010) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5966 ( .A(
        mem_stage_inst_dmem_ram_27__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1011) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5965 ( .A(
        mem_stage_inst_dmem_ram_27__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n1012) );
  NOR2_X0P5A_A12TS mem_stage_inst_dmem_u5964 ( .A(mem_stage_inst_dmem_n218), 
        .B(ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n5951) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5963 ( .A(mem_stage_inst_dmem_n5951), 
        .B(mem_stage_inst_dmem_n165), .C(ex_pipeline_reg_out[24]), .Y(
        mem_stage_inst_dmem_n5698) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5962 ( .A(mem_stage_inst_dmem_n5698), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5969) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5961 ( .A(
        mem_stage_inst_dmem_ram_28__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1013) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5960 ( .A(
        mem_stage_inst_dmem_ram_28__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1014) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5959 ( .A(
        mem_stage_inst_dmem_ram_28__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1015) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5958 ( .A(
        mem_stage_inst_dmem_ram_28__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1016) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5957 ( .A(
        mem_stage_inst_dmem_ram_28__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1017) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5956 ( .A(
        mem_stage_inst_dmem_ram_28__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1018) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5955 ( .A(
        mem_stage_inst_dmem_ram_28__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1019) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5954 ( .A(
        mem_stage_inst_dmem_ram_28__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1020) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5953 ( .A(
        mem_stage_inst_dmem_ram_28__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1021) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5952 ( .A(
        mem_stage_inst_dmem_ram_28__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1022) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5951 ( .A(
        mem_stage_inst_dmem_ram_28__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1023) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5950 ( .A(
        mem_stage_inst_dmem_ram_28__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1024) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5949 ( .A(
        mem_stage_inst_dmem_ram_28__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1025) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5948 ( .A(
        mem_stage_inst_dmem_ram_28__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1026) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5947 ( .A(
        mem_stage_inst_dmem_ram_28__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1027) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5946 ( .A(
        mem_stage_inst_dmem_ram_28__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5969), .Y(mem_stage_inst_dmem_n1028) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5945 ( .A(mem_stage_inst_dmem_n5953), 
        .B(mem_stage_inst_dmem_n166), .C(ex_pipeline_reg_out[24]), .Y(
        mem_stage_inst_dmem_n5696) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5944 ( .A(mem_stage_inst_dmem_n5696), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5968) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5943 ( .A(
        mem_stage_inst_dmem_ram_29__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1029) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5942 ( .A(
        mem_stage_inst_dmem_ram_29__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1030) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5941 ( .A(
        mem_stage_inst_dmem_ram_29__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1031) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5940 ( .A(
        mem_stage_inst_dmem_ram_29__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1032) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5939 ( .A(
        mem_stage_inst_dmem_ram_29__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1033) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5938 ( .A(
        mem_stage_inst_dmem_ram_29__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1034) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5937 ( .A(
        mem_stage_inst_dmem_ram_29__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1035) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5936 ( .A(
        mem_stage_inst_dmem_ram_29__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1036) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5935 ( .A(
        mem_stage_inst_dmem_ram_29__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1037) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5934 ( .A(
        mem_stage_inst_dmem_ram_29__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1038) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5933 ( .A(
        mem_stage_inst_dmem_ram_29__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1039) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5932 ( .A(
        mem_stage_inst_dmem_ram_29__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1040) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5931 ( .A(
        mem_stage_inst_dmem_ram_29__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1041) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5930 ( .A(
        mem_stage_inst_dmem_ram_29__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1042) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5929 ( .A(
        mem_stage_inst_dmem_ram_29__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1043) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5928 ( .A(
        mem_stage_inst_dmem_ram_29__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5968), .Y(mem_stage_inst_dmem_n1044) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5927 ( .A(mem_stage_inst_dmem_n5951), 
        .B(mem_stage_inst_dmem_n164), .C(ex_pipeline_reg_out[24]), .Y(
        mem_stage_inst_dmem_n5694) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5926 ( .A(mem_stage_inst_dmem_n5694), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5967) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5925 ( .A(
        mem_stage_inst_dmem_ram_30__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1045) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5924 ( .A(
        mem_stage_inst_dmem_ram_30__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1046) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5923 ( .A(
        mem_stage_inst_dmem_ram_30__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1047) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5922 ( .A(
        mem_stage_inst_dmem_ram_30__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1048) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5921 ( .A(
        mem_stage_inst_dmem_ram_30__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1049) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5920 ( .A(
        mem_stage_inst_dmem_ram_30__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1050) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5919 ( .A(
        mem_stage_inst_dmem_ram_30__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1051) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5918 ( .A(
        mem_stage_inst_dmem_ram_30__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1052) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5917 ( .A(
        mem_stage_inst_dmem_ram_30__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1053) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5916 ( .A(
        mem_stage_inst_dmem_ram_30__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1054) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5915 ( .A(
        mem_stage_inst_dmem_ram_30__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1055) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5914 ( .A(
        mem_stage_inst_dmem_ram_30__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1056) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5913 ( .A(
        mem_stage_inst_dmem_ram_30__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1057) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5912 ( .A(
        mem_stage_inst_dmem_ram_30__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1058) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5911 ( .A(
        mem_stage_inst_dmem_ram_30__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1059) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5910 ( .A(
        mem_stage_inst_dmem_ram_30__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5967), .Y(mem_stage_inst_dmem_n1060) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5909 ( .A(ex_pipeline_reg_out[23]), 
        .B(mem_stage_inst_dmem_n5953), .C(ex_pipeline_reg_out[24]), .Y(
        mem_stage_inst_dmem_n5691) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5908 ( .A(mem_stage_inst_dmem_n5691), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5966) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5907 ( .A(
        mem_stage_inst_dmem_ram_31__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1061) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5906 ( .A(
        mem_stage_inst_dmem_ram_31__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1062) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5905 ( .A(
        mem_stage_inst_dmem_ram_31__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1063) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5904 ( .A(
        mem_stage_inst_dmem_ram_31__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1064) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5903 ( .A(
        mem_stage_inst_dmem_ram_31__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1065) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5902 ( .A(
        mem_stage_inst_dmem_ram_31__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1066) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5901 ( .A(
        mem_stage_inst_dmem_ram_31__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1067) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5900 ( .A(
        mem_stage_inst_dmem_ram_31__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1068) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5899 ( .A(
        mem_stage_inst_dmem_ram_31__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1069) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5898 ( .A(
        mem_stage_inst_dmem_ram_31__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1070) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5897 ( .A(
        mem_stage_inst_dmem_ram_31__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1071) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5896 ( .A(
        mem_stage_inst_dmem_ram_31__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1072) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5895 ( .A(
        mem_stage_inst_dmem_ram_31__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1073) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5894 ( .A(
        mem_stage_inst_dmem_ram_31__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1074) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5893 ( .A(
        mem_stage_inst_dmem_ram_31__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1075) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5892 ( .A(
        mem_stage_inst_dmem_ram_31__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5966), .Y(mem_stage_inst_dmem_n1076) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5891 ( .A(ex_pipeline_reg_out[27]), 
        .B(mem_stage_inst_dmem_n5965), .Y(mem_stage_inst_dmem_n5750) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5890 ( .A(mem_stage_inst_dmem_n5750), 
        .B(mem_stage_inst_dmem_n5713), .Y(mem_stage_inst_dmem_n5945) );
  NOR2_X0P5A_A12TS mem_stage_inst_dmem_u5889 ( .A(ex_pipeline_reg_out[24]), 
        .B(mem_stage_inst_dmem_n215), .Y(mem_stage_inst_dmem_n5961) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5888 ( .A(mem_stage_inst_dmem_n69), 
        .B(mem_stage_inst_dmem_n167), .C(mem_stage_inst_dmem_n5961), .Y(
        mem_stage_inst_dmem_n5689) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5887 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5964) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5886 ( .A(
        mem_stage_inst_dmem_ram_32__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1077) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5885 ( .A(
        mem_stage_inst_dmem_ram_32__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1078) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5884 ( .A(
        mem_stage_inst_dmem_ram_32__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1079) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5883 ( .A(
        mem_stage_inst_dmem_ram_32__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1080) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5882 ( .A(
        mem_stage_inst_dmem_ram_32__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1081) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5881 ( .A(
        mem_stage_inst_dmem_ram_32__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1082) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5880 ( .A(
        mem_stage_inst_dmem_ram_32__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1083) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5879 ( .A(
        mem_stage_inst_dmem_ram_32__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1084) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5878 ( .A(
        mem_stage_inst_dmem_ram_32__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1085) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5877 ( .A(
        mem_stage_inst_dmem_ram_32__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1086) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5876 ( .A(
        mem_stage_inst_dmem_ram_32__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1087) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5875 ( .A(
        mem_stage_inst_dmem_ram_32__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1088) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5874 ( .A(
        mem_stage_inst_dmem_ram_32__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1089) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5873 ( .A(
        mem_stage_inst_dmem_ram_32__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1090) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5872 ( .A(
        mem_stage_inst_dmem_ram_32__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1091) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5871 ( .A(
        mem_stage_inst_dmem_ram_32__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5964), .Y(mem_stage_inst_dmem_n1092) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5870 ( .A(ex_pipeline_reg_out[22]), 
        .B(mem_stage_inst_dmem_n168), .C(mem_stage_inst_dmem_n5961), .Y(
        mem_stage_inst_dmem_n5687) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5869 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5963) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5868 ( .A(
        mem_stage_inst_dmem_ram_33__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1093) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5867 ( .A(
        mem_stage_inst_dmem_ram_33__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1094) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5866 ( .A(
        mem_stage_inst_dmem_ram_33__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1095) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5865 ( .A(
        mem_stage_inst_dmem_ram_33__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1096) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5864 ( .A(
        mem_stage_inst_dmem_ram_33__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1097) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5863 ( .A(
        mem_stage_inst_dmem_ram_33__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1098) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5862 ( .A(
        mem_stage_inst_dmem_ram_33__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1099) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5861 ( .A(
        mem_stage_inst_dmem_ram_33__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1100) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5860 ( .A(
        mem_stage_inst_dmem_ram_33__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1101) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5859 ( .A(
        mem_stage_inst_dmem_ram_33__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1102) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5858 ( .A(
        mem_stage_inst_dmem_ram_33__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1103) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5857 ( .A(
        mem_stage_inst_dmem_ram_33__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1104) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5856 ( .A(
        mem_stage_inst_dmem_ram_33__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1105) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5855 ( .A(
        mem_stage_inst_dmem_ram_33__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1106) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5854 ( .A(
        mem_stage_inst_dmem_ram_33__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1107) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5853 ( .A(
        mem_stage_inst_dmem_ram_33__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5963), .Y(mem_stage_inst_dmem_n1108) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5852 ( .A(mem_stage_inst_dmem_n164), 
        .B(mem_stage_inst_dmem_n67), .C(mem_stage_inst_dmem_n5961), .Y(
        mem_stage_inst_dmem_n5685) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5851 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5962) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5850 ( .A(
        mem_stage_inst_dmem_ram_34__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1109) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5849 ( .A(
        mem_stage_inst_dmem_ram_34__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1110) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5848 ( .A(
        mem_stage_inst_dmem_ram_34__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1111) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5847 ( .A(
        mem_stage_inst_dmem_ram_34__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1112) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5846 ( .A(
        mem_stage_inst_dmem_ram_34__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1113) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5845 ( .A(
        mem_stage_inst_dmem_ram_34__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1114) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5844 ( .A(
        mem_stage_inst_dmem_ram_34__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1115) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5843 ( .A(
        mem_stage_inst_dmem_ram_34__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1116) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5842 ( .A(
        mem_stage_inst_dmem_ram_34__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1117) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5841 ( .A(
        mem_stage_inst_dmem_ram_34__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1118) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5840 ( .A(
        mem_stage_inst_dmem_ram_34__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1119) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5839 ( .A(
        mem_stage_inst_dmem_ram_34__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1120) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5838 ( .A(
        mem_stage_inst_dmem_ram_34__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1121) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5837 ( .A(
        mem_stage_inst_dmem_ram_34__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1122) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5836 ( .A(
        mem_stage_inst_dmem_ram_34__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1123) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5835 ( .A(
        mem_stage_inst_dmem_ram_34__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5962), .Y(mem_stage_inst_dmem_n1124) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5834 ( .A(mem_stage_inst_dmem_n164), 
        .B(ex_pipeline_reg_out[22]), .C(mem_stage_inst_dmem_n5961), .Y(
        mem_stage_inst_dmem_n5683) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5833 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5960) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5832 ( .A(
        mem_stage_inst_dmem_ram_35__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1125) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5831 ( .A(
        mem_stage_inst_dmem_ram_35__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1126) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5830 ( .A(
        mem_stage_inst_dmem_ram_35__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1127) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5829 ( .A(
        mem_stage_inst_dmem_ram_35__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1128) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5828 ( .A(
        mem_stage_inst_dmem_ram_35__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1129) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5827 ( .A(
        mem_stage_inst_dmem_ram_35__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1130) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5826 ( .A(
        mem_stage_inst_dmem_ram_35__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1131) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5825 ( .A(
        mem_stage_inst_dmem_ram_35__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1132) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5824 ( .A(
        mem_stage_inst_dmem_ram_35__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1133) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5823 ( .A(
        mem_stage_inst_dmem_ram_35__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1134) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5822 ( .A(
        mem_stage_inst_dmem_ram_35__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1135) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5821 ( .A(
        mem_stage_inst_dmem_ram_35__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1136) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5820 ( .A(
        mem_stage_inst_dmem_ram_35__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1137) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5819 ( .A(
        mem_stage_inst_dmem_ram_35__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1138) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5818 ( .A(
        mem_stage_inst_dmem_ram_35__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1139) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5817 ( .A(
        mem_stage_inst_dmem_ram_35__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5960), .Y(mem_stage_inst_dmem_n1140) );
  NOR2_X0P5A_A12TS mem_stage_inst_dmem_u5816 ( .A(mem_stage_inst_dmem_n204), 
        .B(mem_stage_inst_dmem_n209), .Y(mem_stage_inst_dmem_n5956) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5815 ( .A(mem_stage_inst_dmem_n70), 
        .B(mem_stage_inst_dmem_n169), .C(mem_stage_inst_dmem_n5956), .Y(
        mem_stage_inst_dmem_n5681) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5814 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5959) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5813 ( .A(
        mem_stage_inst_dmem_ram_36__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1141) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5812 ( .A(
        mem_stage_inst_dmem_ram_36__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1142) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5811 ( .A(
        mem_stage_inst_dmem_ram_36__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1143) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5810 ( .A(
        mem_stage_inst_dmem_ram_36__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1144) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5809 ( .A(
        mem_stage_inst_dmem_ram_36__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1145) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5808 ( .A(
        mem_stage_inst_dmem_ram_36__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1146) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5807 ( .A(
        mem_stage_inst_dmem_ram_36__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1147) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5806 ( .A(
        mem_stage_inst_dmem_ram_36__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1148) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5805 ( .A(
        mem_stage_inst_dmem_ram_36__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1149) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5804 ( .A(
        mem_stage_inst_dmem_ram_36__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1150) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5803 ( .A(
        mem_stage_inst_dmem_ram_36__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1151) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5802 ( .A(
        mem_stage_inst_dmem_ram_36__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1152) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5801 ( .A(
        mem_stage_inst_dmem_ram_36__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1153) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5800 ( .A(
        mem_stage_inst_dmem_ram_36__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1154) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5799 ( .A(
        mem_stage_inst_dmem_ram_36__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1155) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5798 ( .A(
        mem_stage_inst_dmem_ram_36__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5959), .Y(mem_stage_inst_dmem_n1156) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5797 ( .A(mem_stage_inst_dmem_n40), 
        .B(mem_stage_inst_dmem_n170), .C(mem_stage_inst_dmem_n5956), .Y(
        mem_stage_inst_dmem_n5679) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5796 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5958) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5795 ( .A(
        mem_stage_inst_dmem_ram_37__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1157) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5794 ( .A(
        mem_stage_inst_dmem_ram_37__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1158) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5793 ( .A(
        mem_stage_inst_dmem_ram_37__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1159) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5792 ( .A(
        mem_stage_inst_dmem_ram_37__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1160) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5791 ( .A(
        mem_stage_inst_dmem_ram_37__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1161) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5790 ( .A(
        mem_stage_inst_dmem_ram_37__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1162) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5789 ( .A(
        mem_stage_inst_dmem_ram_37__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1163) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5788 ( .A(
        mem_stage_inst_dmem_ram_37__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1164) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5787 ( .A(
        mem_stage_inst_dmem_ram_37__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1165) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5786 ( .A(
        mem_stage_inst_dmem_ram_37__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1166) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5785 ( .A(
        mem_stage_inst_dmem_ram_37__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1167) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5784 ( .A(
        mem_stage_inst_dmem_ram_37__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1168) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5783 ( .A(
        mem_stage_inst_dmem_ram_37__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1169) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5782 ( .A(
        mem_stage_inst_dmem_ram_37__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1170) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5781 ( .A(
        mem_stage_inst_dmem_ram_37__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1171) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5780 ( .A(
        mem_stage_inst_dmem_ram_37__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5958), .Y(mem_stage_inst_dmem_n1172) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5779 ( .A(mem_stage_inst_dmem_n164), 
        .B(mem_stage_inst_dmem_n68), .C(mem_stage_inst_dmem_n5956), .Y(
        mem_stage_inst_dmem_n5677) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5778 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5957) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5777 ( .A(
        mem_stage_inst_dmem_ram_38__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1173) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5776 ( .A(
        mem_stage_inst_dmem_ram_38__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1174) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5775 ( .A(
        mem_stage_inst_dmem_ram_38__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1175) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5774 ( .A(
        mem_stage_inst_dmem_ram_38__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1176) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5773 ( .A(
        mem_stage_inst_dmem_ram_38__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1177) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5772 ( .A(
        mem_stage_inst_dmem_ram_38__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1178) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5771 ( .A(
        mem_stage_inst_dmem_ram_38__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1179) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5770 ( .A(
        mem_stage_inst_dmem_ram_38__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1180) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5769 ( .A(
        mem_stage_inst_dmem_ram_38__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1181) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5768 ( .A(
        mem_stage_inst_dmem_ram_38__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1182) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5767 ( .A(
        mem_stage_inst_dmem_ram_38__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1183) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5766 ( .A(
        mem_stage_inst_dmem_ram_38__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1184) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5765 ( .A(
        mem_stage_inst_dmem_ram_38__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1185) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5764 ( .A(
        mem_stage_inst_dmem_ram_38__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1186) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5763 ( .A(
        mem_stage_inst_dmem_ram_38__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1187) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5762 ( .A(
        mem_stage_inst_dmem_ram_38__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5957), .Y(mem_stage_inst_dmem_n1188) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5761 ( .A(ex_pipeline_reg_out[23]), 
        .B(ex_pipeline_reg_out[22]), .C(mem_stage_inst_dmem_n5956), .Y(
        mem_stage_inst_dmem_n5675) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5760 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5955) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5759 ( .A(
        mem_stage_inst_dmem_ram_39__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1189) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5758 ( .A(
        mem_stage_inst_dmem_ram_39__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1190) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5757 ( .A(
        mem_stage_inst_dmem_ram_39__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1191) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5756 ( .A(
        mem_stage_inst_dmem_ram_39__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1192) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5755 ( .A(
        mem_stage_inst_dmem_ram_39__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1193) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5754 ( .A(
        mem_stage_inst_dmem_ram_39__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1194) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5753 ( .A(
        mem_stage_inst_dmem_ram_39__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1195) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5752 ( .A(
        mem_stage_inst_dmem_ram_39__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1196) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5751 ( .A(
        mem_stage_inst_dmem_ram_39__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1197) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5750 ( .A(
        mem_stage_inst_dmem_ram_39__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1198) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5749 ( .A(
        mem_stage_inst_dmem_ram_39__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1199) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5748 ( .A(
        mem_stage_inst_dmem_ram_39__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1200) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5747 ( .A(
        mem_stage_inst_dmem_ram_39__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1201) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5746 ( .A(
        mem_stage_inst_dmem_ram_39__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1202) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5745 ( .A(
        mem_stage_inst_dmem_ram_39__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1203) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5744 ( .A(
        mem_stage_inst_dmem_ram_39__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5955), .Y(mem_stage_inst_dmem_n1204) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5743 ( .A(mem_stage_inst_dmem_n171), 
        .B(mem_stage_inst_dmem_n204), .C(mem_stage_inst_dmem_n5951), .Y(
        mem_stage_inst_dmem_n5673) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5742 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5954) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5741 ( .A(
        mem_stage_inst_dmem_ram_40__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1205) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5740 ( .A(
        mem_stage_inst_dmem_ram_40__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1206) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5739 ( .A(
        mem_stage_inst_dmem_ram_40__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1207) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5738 ( .A(
        mem_stage_inst_dmem_ram_40__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1208) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5737 ( .A(
        mem_stage_inst_dmem_ram_40__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1209) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5736 ( .A(
        mem_stage_inst_dmem_ram_40__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1210) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5735 ( .A(
        mem_stage_inst_dmem_ram_40__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1211) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5734 ( .A(
        mem_stage_inst_dmem_ram_40__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1212) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5733 ( .A(
        mem_stage_inst_dmem_ram_40__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1213) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5732 ( .A(
        mem_stage_inst_dmem_ram_40__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1214) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5731 ( .A(
        mem_stage_inst_dmem_ram_40__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1215) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5730 ( .A(
        mem_stage_inst_dmem_ram_40__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1216) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5729 ( .A(
        mem_stage_inst_dmem_ram_40__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1217) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5728 ( .A(
        mem_stage_inst_dmem_ram_40__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1218) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5727 ( .A(
        mem_stage_inst_dmem_ram_40__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1219) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5726 ( .A(
        mem_stage_inst_dmem_ram_40__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5954), .Y(mem_stage_inst_dmem_n1220) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5725 ( .A(mem_stage_inst_dmem_n172), 
        .B(mem_stage_inst_dmem_n204), .C(mem_stage_inst_dmem_n5953), .Y(
        mem_stage_inst_dmem_n5671) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5724 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5952) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5723 ( .A(
        mem_stage_inst_dmem_ram_41__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1221) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5722 ( .A(
        mem_stage_inst_dmem_ram_41__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1222) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5721 ( .A(
        mem_stage_inst_dmem_ram_41__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1223) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5720 ( .A(
        mem_stage_inst_dmem_ram_41__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1224) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5719 ( .A(
        mem_stage_inst_dmem_ram_41__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1225) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5718 ( .A(
        mem_stage_inst_dmem_ram_41__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1226) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5717 ( .A(
        mem_stage_inst_dmem_ram_41__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1227) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5716 ( .A(
        mem_stage_inst_dmem_ram_41__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1228) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5715 ( .A(
        mem_stage_inst_dmem_ram_41__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1229) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5714 ( .A(
        mem_stage_inst_dmem_ram_41__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1230) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5713 ( .A(
        mem_stage_inst_dmem_ram_41__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1231) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5712 ( .A(
        mem_stage_inst_dmem_ram_41__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1232) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5711 ( .A(
        mem_stage_inst_dmem_ram_41__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1233) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5710 ( .A(
        mem_stage_inst_dmem_ram_41__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1234) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5709 ( .A(
        mem_stage_inst_dmem_ram_41__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1235) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5708 ( .A(
        mem_stage_inst_dmem_ram_41__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5952), .Y(mem_stage_inst_dmem_n1236) );
  AND3_X0P5M_A12TS mem_stage_inst_dmem_u5707 ( .A(mem_stage_inst_dmem_n164), 
        .B(mem_stage_inst_dmem_n204), .C(mem_stage_inst_dmem_n5951), .Y(
        mem_stage_inst_dmem_n5668) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5706 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5950) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5705 ( .A(
        mem_stage_inst_dmem_ram_42__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1237) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5704 ( .A(
        mem_stage_inst_dmem_ram_42__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1238) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5703 ( .A(
        mem_stage_inst_dmem_ram_42__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1239) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5702 ( .A(
        mem_stage_inst_dmem_ram_42__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1240) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5701 ( .A(
        mem_stage_inst_dmem_ram_42__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1241) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5700 ( .A(
        mem_stage_inst_dmem_ram_42__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1242) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5699 ( .A(
        mem_stage_inst_dmem_ram_42__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1243) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5698 ( .A(
        mem_stage_inst_dmem_ram_42__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1244) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5697 ( .A(
        mem_stage_inst_dmem_ram_42__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1245) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5696 ( .A(
        mem_stage_inst_dmem_ram_42__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1246) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5695 ( .A(
        mem_stage_inst_dmem_ram_42__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1247) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5694 ( .A(
        mem_stage_inst_dmem_ram_42__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1248) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5693 ( .A(
        mem_stage_inst_dmem_ram_42__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1249) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5692 ( .A(
        mem_stage_inst_dmem_ram_42__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1250) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5691 ( .A(
        mem_stage_inst_dmem_ram_42__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1251) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5690 ( .A(
        mem_stage_inst_dmem_ram_42__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5950), .Y(mem_stage_inst_dmem_n1252) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5689 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5949) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5688 ( .A(
        mem_stage_inst_dmem_ram_43__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1253) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5687 ( .A(
        mem_stage_inst_dmem_ram_43__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1254) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5686 ( .A(
        mem_stage_inst_dmem_ram_43__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1255) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5685 ( .A(
        mem_stage_inst_dmem_ram_43__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1256) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5684 ( .A(
        mem_stage_inst_dmem_ram_43__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1257) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5683 ( .A(
        mem_stage_inst_dmem_ram_43__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1258) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5682 ( .A(
        mem_stage_inst_dmem_ram_43__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1259) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5681 ( .A(
        mem_stage_inst_dmem_ram_43__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1260) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5680 ( .A(
        mem_stage_inst_dmem_ram_43__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1261) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5679 ( .A(
        mem_stage_inst_dmem_ram_43__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1262) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5678 ( .A(
        mem_stage_inst_dmem_ram_43__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1263) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5677 ( .A(
        mem_stage_inst_dmem_ram_43__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1264) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5676 ( .A(
        mem_stage_inst_dmem_ram_43__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1265) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5675 ( .A(
        mem_stage_inst_dmem_ram_43__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1266) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5674 ( .A(
        mem_stage_inst_dmem_ram_43__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1267) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5673 ( .A(
        mem_stage_inst_dmem_ram_43__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5949), .Y(mem_stage_inst_dmem_n1268) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5672 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5948) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5671 ( .A(
        mem_stage_inst_dmem_ram_44__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1269) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5670 ( .A(
        mem_stage_inst_dmem_ram_44__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1270) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5669 ( .A(
        mem_stage_inst_dmem_ram_44__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1271) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5668 ( .A(
        mem_stage_inst_dmem_ram_44__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1272) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5667 ( .A(
        mem_stage_inst_dmem_ram_44__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1273) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5666 ( .A(
        mem_stage_inst_dmem_ram_44__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1274) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5665 ( .A(
        mem_stage_inst_dmem_ram_44__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1275) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5664 ( .A(
        mem_stage_inst_dmem_ram_44__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1276) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5663 ( .A(
        mem_stage_inst_dmem_ram_44__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1277) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5662 ( .A(
        mem_stage_inst_dmem_ram_44__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1278) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5661 ( .A(
        mem_stage_inst_dmem_ram_44__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1279) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5660 ( .A(
        mem_stage_inst_dmem_ram_44__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1280) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5659 ( .A(
        mem_stage_inst_dmem_ram_44__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1281) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5658 ( .A(
        mem_stage_inst_dmem_ram_44__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1282) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5657 ( .A(
        mem_stage_inst_dmem_ram_44__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1283) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5656 ( .A(
        mem_stage_inst_dmem_ram_44__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5948), .Y(mem_stage_inst_dmem_n1284) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5655 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5947) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5654 ( .A(
        mem_stage_inst_dmem_ram_45__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1285) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5653 ( .A(
        mem_stage_inst_dmem_ram_45__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1286) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5652 ( .A(
        mem_stage_inst_dmem_ram_45__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1287) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5651 ( .A(
        mem_stage_inst_dmem_ram_45__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1288) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5650 ( .A(
        mem_stage_inst_dmem_ram_45__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1289) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5649 ( .A(
        mem_stage_inst_dmem_ram_45__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1290) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5648 ( .A(
        mem_stage_inst_dmem_ram_45__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1291) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5647 ( .A(
        mem_stage_inst_dmem_ram_45__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1292) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5646 ( .A(
        mem_stage_inst_dmem_ram_45__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1293) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5645 ( .A(
        mem_stage_inst_dmem_ram_45__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1294) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5644 ( .A(
        mem_stage_inst_dmem_ram_45__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1295) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5643 ( .A(
        mem_stage_inst_dmem_ram_45__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1296) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5642 ( .A(
        mem_stage_inst_dmem_ram_45__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1297) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5641 ( .A(
        mem_stage_inst_dmem_ram_45__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1298) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5640 ( .A(
        mem_stage_inst_dmem_ram_45__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1299) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5639 ( .A(
        mem_stage_inst_dmem_ram_45__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5947), .Y(mem_stage_inst_dmem_n1300) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5638 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5946) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5637 ( .A(
        mem_stage_inst_dmem_ram_46__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1301) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5636 ( .A(
        mem_stage_inst_dmem_ram_46__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1302) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5635 ( .A(
        mem_stage_inst_dmem_ram_46__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1303) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5634 ( .A(
        mem_stage_inst_dmem_ram_46__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1304) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5633 ( .A(
        mem_stage_inst_dmem_ram_46__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1305) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5632 ( .A(
        mem_stage_inst_dmem_ram_46__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1306) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5631 ( .A(
        mem_stage_inst_dmem_ram_46__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1307) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5630 ( .A(
        mem_stage_inst_dmem_ram_46__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1308) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5629 ( .A(
        mem_stage_inst_dmem_ram_46__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1309) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5628 ( .A(
        mem_stage_inst_dmem_ram_46__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1310) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5627 ( .A(
        mem_stage_inst_dmem_ram_46__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1311) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5626 ( .A(
        mem_stage_inst_dmem_ram_46__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1312) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5625 ( .A(
        mem_stage_inst_dmem_ram_46__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1313) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5624 ( .A(
        mem_stage_inst_dmem_ram_46__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1314) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5623 ( .A(
        mem_stage_inst_dmem_ram_46__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1315) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5622 ( .A(
        mem_stage_inst_dmem_ram_46__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5946), .Y(mem_stage_inst_dmem_n1316) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5621 ( .A(mem_stage_inst_dmem_n5945), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5944) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5620 ( .A(
        mem_stage_inst_dmem_ram_47__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1317) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5619 ( .A(
        mem_stage_inst_dmem_ram_47__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1318) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5618 ( .A(
        mem_stage_inst_dmem_ram_47__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1319) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5617 ( .A(
        mem_stage_inst_dmem_ram_47__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1320) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5616 ( .A(
        mem_stage_inst_dmem_ram_47__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1321) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5615 ( .A(
        mem_stage_inst_dmem_ram_47__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1322) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5614 ( .A(
        mem_stage_inst_dmem_ram_47__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1323) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5613 ( .A(
        mem_stage_inst_dmem_ram_47__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1324) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5612 ( .A(
        mem_stage_inst_dmem_ram_47__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1325) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5611 ( .A(
        mem_stage_inst_dmem_ram_47__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1326) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5610 ( .A(
        mem_stage_inst_dmem_ram_47__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1327) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5609 ( .A(
        mem_stage_inst_dmem_ram_47__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1328) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5608 ( .A(
        mem_stage_inst_dmem_ram_47__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1329) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5607 ( .A(
        mem_stage_inst_dmem_ram_47__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1330) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5606 ( .A(
        mem_stage_inst_dmem_ram_47__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1331) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5605 ( .A(
        mem_stage_inst_dmem_ram_47__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5944), .Y(mem_stage_inst_dmem_n1332) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5604 ( .A(ex_pipeline_reg_out[27]), 
        .B(ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5732) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5603 ( .A(mem_stage_inst_dmem_n5732), 
        .B(mem_stage_inst_dmem_n5713), .Y(mem_stage_inst_dmem_n5928) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5602 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5943) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5601 ( .A(
        mem_stage_inst_dmem_ram_48__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1333) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5600 ( .A(
        mem_stage_inst_dmem_ram_48__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1334) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5599 ( .A(
        mem_stage_inst_dmem_ram_48__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1335) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5598 ( .A(
        mem_stage_inst_dmem_ram_48__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1336) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5597 ( .A(
        mem_stage_inst_dmem_ram_48__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1337) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5596 ( .A(
        mem_stage_inst_dmem_ram_48__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1338) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5595 ( .A(
        mem_stage_inst_dmem_ram_48__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1339) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5594 ( .A(
        mem_stage_inst_dmem_ram_48__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1340) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5593 ( .A(
        mem_stage_inst_dmem_ram_48__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1341) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5592 ( .A(
        mem_stage_inst_dmem_ram_48__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1342) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5591 ( .A(
        mem_stage_inst_dmem_ram_48__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1343) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5590 ( .A(
        mem_stage_inst_dmem_ram_48__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1344) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5589 ( .A(
        mem_stage_inst_dmem_ram_48__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1345) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5588 ( .A(
        mem_stage_inst_dmem_ram_48__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1346) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5587 ( .A(
        mem_stage_inst_dmem_ram_48__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1347) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5586 ( .A(
        mem_stage_inst_dmem_ram_48__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5943), .Y(mem_stage_inst_dmem_n1348) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5585 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5942) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5584 ( .A(
        mem_stage_inst_dmem_ram_49__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1349) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5583 ( .A(
        mem_stage_inst_dmem_ram_49__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1350) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5582 ( .A(
        mem_stage_inst_dmem_ram_49__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1351) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5581 ( .A(
        mem_stage_inst_dmem_ram_49__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1352) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5580 ( .A(
        mem_stage_inst_dmem_ram_49__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1353) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5579 ( .A(
        mem_stage_inst_dmem_ram_49__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1354) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5578 ( .A(
        mem_stage_inst_dmem_ram_49__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1355) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5577 ( .A(
        mem_stage_inst_dmem_ram_49__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1356) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5576 ( .A(
        mem_stage_inst_dmem_ram_49__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1357) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5575 ( .A(
        mem_stage_inst_dmem_ram_49__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1358) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5574 ( .A(
        mem_stage_inst_dmem_ram_49__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1359) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5573 ( .A(
        mem_stage_inst_dmem_ram_49__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1360) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5572 ( .A(
        mem_stage_inst_dmem_ram_49__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1361) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5571 ( .A(
        mem_stage_inst_dmem_ram_49__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1362) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5570 ( .A(
        mem_stage_inst_dmem_ram_49__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1363) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5569 ( .A(
        mem_stage_inst_dmem_ram_49__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5942), .Y(mem_stage_inst_dmem_n1364) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5568 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5941) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5567 ( .A(
        mem_stage_inst_dmem_ram_50__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1365) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5566 ( .A(
        mem_stage_inst_dmem_ram_50__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1366) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5565 ( .A(
        mem_stage_inst_dmem_ram_50__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1367) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5564 ( .A(
        mem_stage_inst_dmem_ram_50__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1368) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5563 ( .A(
        mem_stage_inst_dmem_ram_50__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1369) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5562 ( .A(
        mem_stage_inst_dmem_ram_50__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1370) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5561 ( .A(
        mem_stage_inst_dmem_ram_50__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1371) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5560 ( .A(
        mem_stage_inst_dmem_ram_50__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1372) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5559 ( .A(
        mem_stage_inst_dmem_ram_50__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1373) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5558 ( .A(
        mem_stage_inst_dmem_ram_50__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1374) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5557 ( .A(
        mem_stage_inst_dmem_ram_50__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1375) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5556 ( .A(
        mem_stage_inst_dmem_ram_50__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1376) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5555 ( .A(
        mem_stage_inst_dmem_ram_50__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1377) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5554 ( .A(
        mem_stage_inst_dmem_ram_50__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1378) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5553 ( .A(
        mem_stage_inst_dmem_ram_50__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1379) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5552 ( .A(
        mem_stage_inst_dmem_ram_50__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5941), .Y(mem_stage_inst_dmem_n1380) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5551 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5940) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5550 ( .A(
        mem_stage_inst_dmem_ram_51__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1381) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5549 ( .A(
        mem_stage_inst_dmem_ram_51__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1382) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5548 ( .A(
        mem_stage_inst_dmem_ram_51__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1383) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5547 ( .A(
        mem_stage_inst_dmem_ram_51__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1384) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5546 ( .A(
        mem_stage_inst_dmem_ram_51__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1385) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5545 ( .A(
        mem_stage_inst_dmem_ram_51__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1386) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5544 ( .A(
        mem_stage_inst_dmem_ram_51__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1387) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5543 ( .A(
        mem_stage_inst_dmem_ram_51__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1388) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5542 ( .A(
        mem_stage_inst_dmem_ram_51__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1389) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5541 ( .A(
        mem_stage_inst_dmem_ram_51__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1390) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5540 ( .A(
        mem_stage_inst_dmem_ram_51__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1391) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5539 ( .A(
        mem_stage_inst_dmem_ram_51__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1392) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5538 ( .A(
        mem_stage_inst_dmem_ram_51__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1393) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5537 ( .A(
        mem_stage_inst_dmem_ram_51__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1394) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5536 ( .A(
        mem_stage_inst_dmem_ram_51__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1395) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5535 ( .A(
        mem_stage_inst_dmem_ram_51__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5940), .Y(mem_stage_inst_dmem_n1396) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5534 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5939) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5533 ( .A(
        mem_stage_inst_dmem_ram_52__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1397) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5532 ( .A(
        mem_stage_inst_dmem_ram_52__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1398) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5531 ( .A(
        mem_stage_inst_dmem_ram_52__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1399) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5530 ( .A(
        mem_stage_inst_dmem_ram_52__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1400) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5529 ( .A(
        mem_stage_inst_dmem_ram_52__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1401) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5528 ( .A(
        mem_stage_inst_dmem_ram_52__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1402) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5527 ( .A(
        mem_stage_inst_dmem_ram_52__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1403) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5526 ( .A(
        mem_stage_inst_dmem_ram_52__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1404) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5525 ( .A(
        mem_stage_inst_dmem_ram_52__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1405) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5524 ( .A(
        mem_stage_inst_dmem_ram_52__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1406) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5523 ( .A(
        mem_stage_inst_dmem_ram_52__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1407) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5522 ( .A(
        mem_stage_inst_dmem_ram_52__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1408) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5521 ( .A(
        mem_stage_inst_dmem_ram_52__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1409) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5520 ( .A(
        mem_stage_inst_dmem_ram_52__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1410) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5519 ( .A(
        mem_stage_inst_dmem_ram_52__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1411) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5518 ( .A(
        mem_stage_inst_dmem_ram_52__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5939), .Y(mem_stage_inst_dmem_n1412) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5517 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5938) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5516 ( .A(
        mem_stage_inst_dmem_ram_53__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1413) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5515 ( .A(
        mem_stage_inst_dmem_ram_53__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1414) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5514 ( .A(
        mem_stage_inst_dmem_ram_53__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1415) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5513 ( .A(
        mem_stage_inst_dmem_ram_53__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1416) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5512 ( .A(
        mem_stage_inst_dmem_ram_53__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1417) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5511 ( .A(
        mem_stage_inst_dmem_ram_53__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1418) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5510 ( .A(
        mem_stage_inst_dmem_ram_53__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1419) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5509 ( .A(
        mem_stage_inst_dmem_ram_53__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1420) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5508 ( .A(
        mem_stage_inst_dmem_ram_53__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1421) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5507 ( .A(
        mem_stage_inst_dmem_ram_53__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1422) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5506 ( .A(
        mem_stage_inst_dmem_ram_53__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1423) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5505 ( .A(
        mem_stage_inst_dmem_ram_53__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1424) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5504 ( .A(
        mem_stage_inst_dmem_ram_53__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1425) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5503 ( .A(
        mem_stage_inst_dmem_ram_53__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1426) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5502 ( .A(
        mem_stage_inst_dmem_ram_53__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1427) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5501 ( .A(
        mem_stage_inst_dmem_ram_53__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5938), .Y(mem_stage_inst_dmem_n1428) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5500 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5937) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5499 ( .A(
        mem_stage_inst_dmem_ram_54__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1429) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5498 ( .A(
        mem_stage_inst_dmem_ram_54__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1430) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5497 ( .A(
        mem_stage_inst_dmem_ram_54__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1431) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5496 ( .A(
        mem_stage_inst_dmem_ram_54__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1432) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5495 ( .A(
        mem_stage_inst_dmem_ram_54__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1433) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5494 ( .A(
        mem_stage_inst_dmem_ram_54__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1434) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5493 ( .A(
        mem_stage_inst_dmem_ram_54__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1435) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5492 ( .A(
        mem_stage_inst_dmem_ram_54__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1436) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5491 ( .A(
        mem_stage_inst_dmem_ram_54__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1437) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5490 ( .A(
        mem_stage_inst_dmem_ram_54__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1438) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5489 ( .A(
        mem_stage_inst_dmem_ram_54__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1439) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5488 ( .A(
        mem_stage_inst_dmem_ram_54__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1440) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5487 ( .A(
        mem_stage_inst_dmem_ram_54__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1441) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5486 ( .A(
        mem_stage_inst_dmem_ram_54__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1442) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5485 ( .A(
        mem_stage_inst_dmem_ram_54__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1443) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5484 ( .A(
        mem_stage_inst_dmem_ram_54__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5937), .Y(mem_stage_inst_dmem_n1444) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5483 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5936) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5482 ( .A(
        mem_stage_inst_dmem_ram_55__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1445) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5481 ( .A(
        mem_stage_inst_dmem_ram_55__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1446) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5480 ( .A(
        mem_stage_inst_dmem_ram_55__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1447) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5479 ( .A(
        mem_stage_inst_dmem_ram_55__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1448) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5478 ( .A(
        mem_stage_inst_dmem_ram_55__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1449) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5477 ( .A(
        mem_stage_inst_dmem_ram_55__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1450) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5476 ( .A(
        mem_stage_inst_dmem_ram_55__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1451) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5475 ( .A(
        mem_stage_inst_dmem_ram_55__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1452) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5474 ( .A(
        mem_stage_inst_dmem_ram_55__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1453) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5473 ( .A(
        mem_stage_inst_dmem_ram_55__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1454) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5472 ( .A(
        mem_stage_inst_dmem_ram_55__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1455) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5471 ( .A(
        mem_stage_inst_dmem_ram_55__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1456) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5470 ( .A(
        mem_stage_inst_dmem_ram_55__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1457) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5469 ( .A(
        mem_stage_inst_dmem_ram_55__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1458) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5468 ( .A(
        mem_stage_inst_dmem_ram_55__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1459) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5467 ( .A(
        mem_stage_inst_dmem_ram_55__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5936), .Y(mem_stage_inst_dmem_n1460) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5466 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5935) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5465 ( .A(
        mem_stage_inst_dmem_ram_56__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1461) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5464 ( .A(
        mem_stage_inst_dmem_ram_56__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1462) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5463 ( .A(
        mem_stage_inst_dmem_ram_56__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1463) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5462 ( .A(
        mem_stage_inst_dmem_ram_56__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1464) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5461 ( .A(
        mem_stage_inst_dmem_ram_56__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1465) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5460 ( .A(
        mem_stage_inst_dmem_ram_56__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1466) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5459 ( .A(
        mem_stage_inst_dmem_ram_56__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1467) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5458 ( .A(
        mem_stage_inst_dmem_ram_56__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1468) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5457 ( .A(
        mem_stage_inst_dmem_ram_56__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1469) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5456 ( .A(
        mem_stage_inst_dmem_ram_56__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1470) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5455 ( .A(
        mem_stage_inst_dmem_ram_56__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1471) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5454 ( .A(
        mem_stage_inst_dmem_ram_56__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1472) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5453 ( .A(
        mem_stage_inst_dmem_ram_56__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1473) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5452 ( .A(
        mem_stage_inst_dmem_ram_56__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1474) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5451 ( .A(
        mem_stage_inst_dmem_ram_56__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1475) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5450 ( .A(
        mem_stage_inst_dmem_ram_56__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5935), .Y(mem_stage_inst_dmem_n1476) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5449 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5934) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5448 ( .A(
        mem_stage_inst_dmem_ram_57__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1477) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5447 ( .A(
        mem_stage_inst_dmem_ram_57__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1478) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5446 ( .A(
        mem_stage_inst_dmem_ram_57__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1479) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5445 ( .A(
        mem_stage_inst_dmem_ram_57__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1480) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5444 ( .A(
        mem_stage_inst_dmem_ram_57__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1481) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5443 ( .A(
        mem_stage_inst_dmem_ram_57__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1482) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5442 ( .A(
        mem_stage_inst_dmem_ram_57__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1483) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5441 ( .A(
        mem_stage_inst_dmem_ram_57__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1484) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5440 ( .A(
        mem_stage_inst_dmem_ram_57__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1485) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5439 ( .A(
        mem_stage_inst_dmem_ram_57__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1486) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5438 ( .A(
        mem_stage_inst_dmem_ram_57__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1487) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5437 ( .A(
        mem_stage_inst_dmem_ram_57__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1488) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5436 ( .A(
        mem_stage_inst_dmem_ram_57__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1489) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5435 ( .A(
        mem_stage_inst_dmem_ram_57__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1490) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5434 ( .A(
        mem_stage_inst_dmem_ram_57__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1491) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5433 ( .A(
        mem_stage_inst_dmem_ram_57__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5934), .Y(mem_stage_inst_dmem_n1492) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5432 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5933) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5431 ( .A(
        mem_stage_inst_dmem_ram_58__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1493) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5430 ( .A(
        mem_stage_inst_dmem_ram_58__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1494) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5429 ( .A(
        mem_stage_inst_dmem_ram_58__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1495) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5428 ( .A(
        mem_stage_inst_dmem_ram_58__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1496) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5427 ( .A(
        mem_stage_inst_dmem_ram_58__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1497) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5426 ( .A(
        mem_stage_inst_dmem_ram_58__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1498) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5425 ( .A(
        mem_stage_inst_dmem_ram_58__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1499) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5424 ( .A(
        mem_stage_inst_dmem_ram_58__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1500) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5423 ( .A(
        mem_stage_inst_dmem_ram_58__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1501) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5422 ( .A(
        mem_stage_inst_dmem_ram_58__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1502) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5421 ( .A(
        mem_stage_inst_dmem_ram_58__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1503) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5420 ( .A(
        mem_stage_inst_dmem_ram_58__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1504) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5419 ( .A(
        mem_stage_inst_dmem_ram_58__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1505) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5418 ( .A(
        mem_stage_inst_dmem_ram_58__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1506) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5417 ( .A(
        mem_stage_inst_dmem_ram_58__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1507) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5416 ( .A(
        mem_stage_inst_dmem_ram_58__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5933), .Y(mem_stage_inst_dmem_n1508) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5415 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5932) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5414 ( .A(
        mem_stage_inst_dmem_ram_59__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1509) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5413 ( .A(
        mem_stage_inst_dmem_ram_59__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1510) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5412 ( .A(
        mem_stage_inst_dmem_ram_59__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1511) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5411 ( .A(
        mem_stage_inst_dmem_ram_59__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1512) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5410 ( .A(
        mem_stage_inst_dmem_ram_59__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1513) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5409 ( .A(
        mem_stage_inst_dmem_ram_59__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1514) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5408 ( .A(
        mem_stage_inst_dmem_ram_59__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1515) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5407 ( .A(
        mem_stage_inst_dmem_ram_59__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1516) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5406 ( .A(
        mem_stage_inst_dmem_ram_59__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1517) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5405 ( .A(
        mem_stage_inst_dmem_ram_59__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1518) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5404 ( .A(
        mem_stage_inst_dmem_ram_59__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1519) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5403 ( .A(
        mem_stage_inst_dmem_ram_59__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1520) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5402 ( .A(
        mem_stage_inst_dmem_ram_59__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1521) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5401 ( .A(
        mem_stage_inst_dmem_ram_59__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1522) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5400 ( .A(
        mem_stage_inst_dmem_ram_59__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1523) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5399 ( .A(
        mem_stage_inst_dmem_ram_59__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5932), .Y(mem_stage_inst_dmem_n1524) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5398 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5931) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5397 ( .A(
        mem_stage_inst_dmem_ram_60__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1525) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5396 ( .A(
        mem_stage_inst_dmem_ram_60__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1526) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5395 ( .A(
        mem_stage_inst_dmem_ram_60__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1527) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5394 ( .A(
        mem_stage_inst_dmem_ram_60__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1528) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5393 ( .A(
        mem_stage_inst_dmem_ram_60__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1529) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5392 ( .A(
        mem_stage_inst_dmem_ram_60__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1530) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5391 ( .A(
        mem_stage_inst_dmem_ram_60__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1531) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5390 ( .A(
        mem_stage_inst_dmem_ram_60__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1532) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5389 ( .A(
        mem_stage_inst_dmem_ram_60__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1533) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5388 ( .A(
        mem_stage_inst_dmem_ram_60__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1534) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5387 ( .A(
        mem_stage_inst_dmem_ram_60__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1535) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5386 ( .A(
        mem_stage_inst_dmem_ram_60__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1536) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5385 ( .A(
        mem_stage_inst_dmem_ram_60__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1537) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5384 ( .A(
        mem_stage_inst_dmem_ram_60__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1538) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5383 ( .A(
        mem_stage_inst_dmem_ram_60__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1539) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5382 ( .A(
        mem_stage_inst_dmem_ram_60__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5931), .Y(mem_stage_inst_dmem_n1540) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5381 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5930) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5380 ( .A(
        mem_stage_inst_dmem_ram_61__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1541) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5379 ( .A(
        mem_stage_inst_dmem_ram_61__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1542) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5378 ( .A(
        mem_stage_inst_dmem_ram_61__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1543) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5377 ( .A(
        mem_stage_inst_dmem_ram_61__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1544) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5376 ( .A(
        mem_stage_inst_dmem_ram_61__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1545) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5375 ( .A(
        mem_stage_inst_dmem_ram_61__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1546) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5374 ( .A(
        mem_stage_inst_dmem_ram_61__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1547) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5373 ( .A(
        mem_stage_inst_dmem_ram_61__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1548) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5372 ( .A(
        mem_stage_inst_dmem_ram_61__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1549) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5371 ( .A(
        mem_stage_inst_dmem_ram_61__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1550) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5370 ( .A(
        mem_stage_inst_dmem_ram_61__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1551) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5369 ( .A(
        mem_stage_inst_dmem_ram_61__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1552) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5368 ( .A(
        mem_stage_inst_dmem_ram_61__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1553) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5367 ( .A(
        mem_stage_inst_dmem_ram_61__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1554) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5366 ( .A(
        mem_stage_inst_dmem_ram_61__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1555) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5365 ( .A(
        mem_stage_inst_dmem_ram_61__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5930), .Y(mem_stage_inst_dmem_n1556) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5364 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5929) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5363 ( .A(
        mem_stage_inst_dmem_ram_62__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1557) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5362 ( .A(
        mem_stage_inst_dmem_ram_62__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1558) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5361 ( .A(
        mem_stage_inst_dmem_ram_62__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1559) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5360 ( .A(
        mem_stage_inst_dmem_ram_62__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1560) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5359 ( .A(
        mem_stage_inst_dmem_ram_62__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1561) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5358 ( .A(
        mem_stage_inst_dmem_ram_62__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1562) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5357 ( .A(
        mem_stage_inst_dmem_ram_62__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1563) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5356 ( .A(
        mem_stage_inst_dmem_ram_62__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1564) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5355 ( .A(
        mem_stage_inst_dmem_ram_62__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1565) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5354 ( .A(
        mem_stage_inst_dmem_ram_62__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1566) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5353 ( .A(
        mem_stage_inst_dmem_ram_62__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1567) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5352 ( .A(
        mem_stage_inst_dmem_ram_62__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1568) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5351 ( .A(
        mem_stage_inst_dmem_ram_62__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1569) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5350 ( .A(
        mem_stage_inst_dmem_ram_62__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1570) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5349 ( .A(
        mem_stage_inst_dmem_ram_62__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1571) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5348 ( .A(
        mem_stage_inst_dmem_ram_62__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5929), .Y(mem_stage_inst_dmem_n1572) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5347 ( .A(mem_stage_inst_dmem_n5928), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5927) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5346 ( .A(
        mem_stage_inst_dmem_ram_63__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1573) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5345 ( .A(
        mem_stage_inst_dmem_ram_63__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1574) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5344 ( .A(
        mem_stage_inst_dmem_ram_63__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1575) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5343 ( .A(
        mem_stage_inst_dmem_ram_63__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1576) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5342 ( .A(
        mem_stage_inst_dmem_ram_63__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1577) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5341 ( .A(
        mem_stage_inst_dmem_ram_63__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1578) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5340 ( .A(
        mem_stage_inst_dmem_ram_63__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1579) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5339 ( .A(
        mem_stage_inst_dmem_ram_63__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1580) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5338 ( .A(
        mem_stage_inst_dmem_ram_63__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1581) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5337 ( .A(
        mem_stage_inst_dmem_ram_63__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1582) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5336 ( .A(
        mem_stage_inst_dmem_ram_63__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1583) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5335 ( .A(
        mem_stage_inst_dmem_ram_63__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1584) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5334 ( .A(
        mem_stage_inst_dmem_ram_63__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1585) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5333 ( .A(
        mem_stage_inst_dmem_ram_63__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1586) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5332 ( .A(
        mem_stage_inst_dmem_ram_63__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1587) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5331 ( .A(
        mem_stage_inst_dmem_ram_63__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5927), .Y(mem_stage_inst_dmem_n1588) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5330 ( .A(mem_stage_inst_dmem_n5926), 
        .B(ex_pipeline_reg_out[28]), .Y(mem_stage_inst_dmem_n5874) );
  NOR2_X0P5A_A12TS mem_stage_inst_dmem_u5329 ( .A(ex_pipeline_reg_out[26]), 
        .B(ex_pipeline_reg_out[27]), .Y(mem_stage_inst_dmem_n5712) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5328 ( .A(mem_stage_inst_dmem_n5874), 
        .B(mem_stage_inst_dmem_n5712), .Y(mem_stage_inst_dmem_n5910) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5327 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5925) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5326 ( .A(
        mem_stage_inst_dmem_ram_64__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1589) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5325 ( .A(
        mem_stage_inst_dmem_ram_64__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1590) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5324 ( .A(
        mem_stage_inst_dmem_ram_64__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1591) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5323 ( .A(
        mem_stage_inst_dmem_ram_64__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1592) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5322 ( .A(
        mem_stage_inst_dmem_ram_64__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1593) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5321 ( .A(
        mem_stage_inst_dmem_ram_64__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1594) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5320 ( .A(
        mem_stage_inst_dmem_ram_64__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1595) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5319 ( .A(
        mem_stage_inst_dmem_ram_64__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1596) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5318 ( .A(
        mem_stage_inst_dmem_ram_64__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1597) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5317 ( .A(
        mem_stage_inst_dmem_ram_64__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1598) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5316 ( .A(
        mem_stage_inst_dmem_ram_64__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1599) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5315 ( .A(
        mem_stage_inst_dmem_ram_64__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1600) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5314 ( .A(
        mem_stage_inst_dmem_ram_64__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1601) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5313 ( .A(
        mem_stage_inst_dmem_ram_64__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1602) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5312 ( .A(
        mem_stage_inst_dmem_ram_64__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1603) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5311 ( .A(
        mem_stage_inst_dmem_ram_64__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5925), .Y(mem_stage_inst_dmem_n1604) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5310 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5924) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5309 ( .A(
        mem_stage_inst_dmem_ram_65__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1605) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5308 ( .A(
        mem_stage_inst_dmem_ram_65__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1606) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5307 ( .A(
        mem_stage_inst_dmem_ram_65__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1607) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5306 ( .A(
        mem_stage_inst_dmem_ram_65__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1608) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5305 ( .A(
        mem_stage_inst_dmem_ram_65__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1609) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5304 ( .A(
        mem_stage_inst_dmem_ram_65__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1610) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5303 ( .A(
        mem_stage_inst_dmem_ram_65__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1611) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5302 ( .A(
        mem_stage_inst_dmem_ram_65__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1612) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5301 ( .A(
        mem_stage_inst_dmem_ram_65__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1613) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5300 ( .A(
        mem_stage_inst_dmem_ram_65__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1614) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5299 ( .A(
        mem_stage_inst_dmem_ram_65__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1615) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5298 ( .A(
        mem_stage_inst_dmem_ram_65__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1616) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5297 ( .A(
        mem_stage_inst_dmem_ram_65__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1617) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5296 ( .A(
        mem_stage_inst_dmem_ram_65__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1618) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5295 ( .A(
        mem_stage_inst_dmem_ram_65__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1619) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5294 ( .A(
        mem_stage_inst_dmem_ram_65__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5924), .Y(mem_stage_inst_dmem_n1620) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5293 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5923) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5292 ( .A(
        mem_stage_inst_dmem_ram_66__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1621) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5291 ( .A(
        mem_stage_inst_dmem_ram_66__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1622) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5290 ( .A(
        mem_stage_inst_dmem_ram_66__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1623) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5289 ( .A(
        mem_stage_inst_dmem_ram_66__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1624) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5288 ( .A(
        mem_stage_inst_dmem_ram_66__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1625) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5287 ( .A(
        mem_stage_inst_dmem_ram_66__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1626) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5286 ( .A(
        mem_stage_inst_dmem_ram_66__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1627) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5285 ( .A(
        mem_stage_inst_dmem_ram_66__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1628) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5284 ( .A(
        mem_stage_inst_dmem_ram_66__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1629) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5283 ( .A(
        mem_stage_inst_dmem_ram_66__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1630) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5282 ( .A(
        mem_stage_inst_dmem_ram_66__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1631) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5281 ( .A(
        mem_stage_inst_dmem_ram_66__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1632) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5280 ( .A(
        mem_stage_inst_dmem_ram_66__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1633) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5279 ( .A(
        mem_stage_inst_dmem_ram_66__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1634) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5278 ( .A(
        mem_stage_inst_dmem_ram_66__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1635) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5277 ( .A(
        mem_stage_inst_dmem_ram_66__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5923), .Y(mem_stage_inst_dmem_n1636) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5276 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5922) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5275 ( .A(
        mem_stage_inst_dmem_ram_67__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1637) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5274 ( .A(
        mem_stage_inst_dmem_ram_67__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1638) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5273 ( .A(
        mem_stage_inst_dmem_ram_67__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1639) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5272 ( .A(
        mem_stage_inst_dmem_ram_67__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1640) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5271 ( .A(
        mem_stage_inst_dmem_ram_67__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1641) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5270 ( .A(
        mem_stage_inst_dmem_ram_67__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1642) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5269 ( .A(
        mem_stage_inst_dmem_ram_67__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1643) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5268 ( .A(
        mem_stage_inst_dmem_ram_67__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1644) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5267 ( .A(
        mem_stage_inst_dmem_ram_67__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1645) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5266 ( .A(
        mem_stage_inst_dmem_ram_67__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1646) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5265 ( .A(
        mem_stage_inst_dmem_ram_67__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1647) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5264 ( .A(
        mem_stage_inst_dmem_ram_67__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1648) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5263 ( .A(
        mem_stage_inst_dmem_ram_67__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1649) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5262 ( .A(
        mem_stage_inst_dmem_ram_67__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1650) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5261 ( .A(
        mem_stage_inst_dmem_ram_67__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1651) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5260 ( .A(
        mem_stage_inst_dmem_ram_67__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5922), .Y(mem_stage_inst_dmem_n1652) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5259 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5921) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5258 ( .A(
        mem_stage_inst_dmem_ram_68__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1653) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5257 ( .A(
        mem_stage_inst_dmem_ram_68__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1654) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5256 ( .A(
        mem_stage_inst_dmem_ram_68__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1655) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5255 ( .A(
        mem_stage_inst_dmem_ram_68__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1656) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5254 ( .A(
        mem_stage_inst_dmem_ram_68__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1657) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5253 ( .A(
        mem_stage_inst_dmem_ram_68__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1658) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5252 ( .A(
        mem_stage_inst_dmem_ram_68__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1659) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5251 ( .A(
        mem_stage_inst_dmem_ram_68__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1660) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5250 ( .A(
        mem_stage_inst_dmem_ram_68__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1661) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5249 ( .A(
        mem_stage_inst_dmem_ram_68__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1662) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5248 ( .A(
        mem_stage_inst_dmem_ram_68__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1663) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5247 ( .A(
        mem_stage_inst_dmem_ram_68__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1664) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5246 ( .A(
        mem_stage_inst_dmem_ram_68__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1665) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5245 ( .A(
        mem_stage_inst_dmem_ram_68__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1666) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5244 ( .A(
        mem_stage_inst_dmem_ram_68__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1667) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5243 ( .A(
        mem_stage_inst_dmem_ram_68__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5921), .Y(mem_stage_inst_dmem_n1668) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5242 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5920) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5241 ( .A(
        mem_stage_inst_dmem_ram_69__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1669) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5240 ( .A(
        mem_stage_inst_dmem_ram_69__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1670) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5239 ( .A(
        mem_stage_inst_dmem_ram_69__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1671) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5238 ( .A(
        mem_stage_inst_dmem_ram_69__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1672) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5237 ( .A(
        mem_stage_inst_dmem_ram_69__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1673) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5236 ( .A(
        mem_stage_inst_dmem_ram_69__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1674) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5235 ( .A(
        mem_stage_inst_dmem_ram_69__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1675) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5234 ( .A(
        mem_stage_inst_dmem_ram_69__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1676) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5233 ( .A(
        mem_stage_inst_dmem_ram_69__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1677) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5232 ( .A(
        mem_stage_inst_dmem_ram_69__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1678) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5231 ( .A(
        mem_stage_inst_dmem_ram_69__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1679) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5230 ( .A(
        mem_stage_inst_dmem_ram_69__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1680) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5229 ( .A(
        mem_stage_inst_dmem_ram_69__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1681) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5228 ( .A(
        mem_stage_inst_dmem_ram_69__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1682) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5227 ( .A(
        mem_stage_inst_dmem_ram_69__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1683) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5226 ( .A(
        mem_stage_inst_dmem_ram_69__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5920), .Y(mem_stage_inst_dmem_n1684) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5225 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5919) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5224 ( .A(
        mem_stage_inst_dmem_ram_70__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1685) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5223 ( .A(
        mem_stage_inst_dmem_ram_70__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1686) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5222 ( .A(
        mem_stage_inst_dmem_ram_70__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1687) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5221 ( .A(
        mem_stage_inst_dmem_ram_70__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1688) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5220 ( .A(
        mem_stage_inst_dmem_ram_70__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1689) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5219 ( .A(
        mem_stage_inst_dmem_ram_70__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1690) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5218 ( .A(
        mem_stage_inst_dmem_ram_70__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1691) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5217 ( .A(
        mem_stage_inst_dmem_ram_70__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1692) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5216 ( .A(
        mem_stage_inst_dmem_ram_70__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1693) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5215 ( .A(
        mem_stage_inst_dmem_ram_70__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1694) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5214 ( .A(
        mem_stage_inst_dmem_ram_70__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1695) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5213 ( .A(
        mem_stage_inst_dmem_ram_70__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1696) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5212 ( .A(
        mem_stage_inst_dmem_ram_70__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1697) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5211 ( .A(
        mem_stage_inst_dmem_ram_70__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1698) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5210 ( .A(
        mem_stage_inst_dmem_ram_70__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1699) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5209 ( .A(
        mem_stage_inst_dmem_ram_70__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5919), .Y(mem_stage_inst_dmem_n1700) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5208 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5918) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5207 ( .A(
        mem_stage_inst_dmem_ram_71__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1701) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5206 ( .A(
        mem_stage_inst_dmem_ram_71__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1702) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5205 ( .A(
        mem_stage_inst_dmem_ram_71__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1703) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5204 ( .A(
        mem_stage_inst_dmem_ram_71__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1704) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5203 ( .A(
        mem_stage_inst_dmem_ram_71__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1705) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5202 ( .A(
        mem_stage_inst_dmem_ram_71__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1706) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5201 ( .A(
        mem_stage_inst_dmem_ram_71__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1707) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5200 ( .A(
        mem_stage_inst_dmem_ram_71__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1708) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5199 ( .A(
        mem_stage_inst_dmem_ram_71__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1709) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5198 ( .A(
        mem_stage_inst_dmem_ram_71__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1710) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5197 ( .A(
        mem_stage_inst_dmem_ram_71__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1711) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5196 ( .A(
        mem_stage_inst_dmem_ram_71__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1712) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5195 ( .A(
        mem_stage_inst_dmem_ram_71__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1713) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5194 ( .A(
        mem_stage_inst_dmem_ram_71__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1714) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5193 ( .A(
        mem_stage_inst_dmem_ram_71__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1715) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5192 ( .A(
        mem_stage_inst_dmem_ram_71__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5918), .Y(mem_stage_inst_dmem_n1716) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5191 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5917) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5190 ( .A(
        mem_stage_inst_dmem_ram_72__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1717) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5189 ( .A(
        mem_stage_inst_dmem_ram_72__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1718) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5188 ( .A(
        mem_stage_inst_dmem_ram_72__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1719) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5187 ( .A(
        mem_stage_inst_dmem_ram_72__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1720) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5186 ( .A(
        mem_stage_inst_dmem_ram_72__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1721) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5185 ( .A(
        mem_stage_inst_dmem_ram_72__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1722) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5184 ( .A(
        mem_stage_inst_dmem_ram_72__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1723) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5183 ( .A(
        mem_stage_inst_dmem_ram_72__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1724) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5182 ( .A(
        mem_stage_inst_dmem_ram_72__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1725) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5181 ( .A(
        mem_stage_inst_dmem_ram_72__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1726) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5180 ( .A(
        mem_stage_inst_dmem_ram_72__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1727) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5179 ( .A(
        mem_stage_inst_dmem_ram_72__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1728) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5178 ( .A(
        mem_stage_inst_dmem_ram_72__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1729) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5177 ( .A(
        mem_stage_inst_dmem_ram_72__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1730) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5176 ( .A(
        mem_stage_inst_dmem_ram_72__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1731) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5175 ( .A(
        mem_stage_inst_dmem_ram_72__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5917), .Y(mem_stage_inst_dmem_n1732) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5174 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5916) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5173 ( .A(
        mem_stage_inst_dmem_ram_73__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1733) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5172 ( .A(
        mem_stage_inst_dmem_ram_73__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1734) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5171 ( .A(
        mem_stage_inst_dmem_ram_73__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1735) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5170 ( .A(
        mem_stage_inst_dmem_ram_73__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1736) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5169 ( .A(
        mem_stage_inst_dmem_ram_73__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1737) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5168 ( .A(
        mem_stage_inst_dmem_ram_73__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1738) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5167 ( .A(
        mem_stage_inst_dmem_ram_73__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1739) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5166 ( .A(
        mem_stage_inst_dmem_ram_73__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1740) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5165 ( .A(
        mem_stage_inst_dmem_ram_73__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1741) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5164 ( .A(
        mem_stage_inst_dmem_ram_73__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1742) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5163 ( .A(
        mem_stage_inst_dmem_ram_73__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1743) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5162 ( .A(
        mem_stage_inst_dmem_ram_73__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1744) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5161 ( .A(
        mem_stage_inst_dmem_ram_73__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1745) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5160 ( .A(
        mem_stage_inst_dmem_ram_73__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1746) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5159 ( .A(
        mem_stage_inst_dmem_ram_73__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1747) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5158 ( .A(
        mem_stage_inst_dmem_ram_73__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5916), .Y(mem_stage_inst_dmem_n1748) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5157 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5915) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5156 ( .A(
        mem_stage_inst_dmem_ram_74__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1749) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5155 ( .A(
        mem_stage_inst_dmem_ram_74__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1750) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5154 ( .A(
        mem_stage_inst_dmem_ram_74__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1751) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5153 ( .A(
        mem_stage_inst_dmem_ram_74__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1752) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5152 ( .A(
        mem_stage_inst_dmem_ram_74__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1753) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5151 ( .A(
        mem_stage_inst_dmem_ram_74__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1754) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5150 ( .A(
        mem_stage_inst_dmem_ram_74__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1755) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5149 ( .A(
        mem_stage_inst_dmem_ram_74__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1756) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5148 ( .A(
        mem_stage_inst_dmem_ram_74__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1757) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5147 ( .A(
        mem_stage_inst_dmem_ram_74__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1758) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5146 ( .A(
        mem_stage_inst_dmem_ram_74__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1759) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5145 ( .A(
        mem_stage_inst_dmem_ram_74__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1760) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5144 ( .A(
        mem_stage_inst_dmem_ram_74__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1761) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5143 ( .A(
        mem_stage_inst_dmem_ram_74__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1762) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5142 ( .A(
        mem_stage_inst_dmem_ram_74__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1763) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5141 ( .A(
        mem_stage_inst_dmem_ram_74__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5915), .Y(mem_stage_inst_dmem_n1764) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5140 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5914) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5139 ( .A(
        mem_stage_inst_dmem_ram_75__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1765) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5138 ( .A(
        mem_stage_inst_dmem_ram_75__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1766) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5137 ( .A(
        mem_stage_inst_dmem_ram_75__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1767) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5136 ( .A(
        mem_stage_inst_dmem_ram_75__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1768) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5135 ( .A(
        mem_stage_inst_dmem_ram_75__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1769) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5134 ( .A(
        mem_stage_inst_dmem_ram_75__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1770) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5133 ( .A(
        mem_stage_inst_dmem_ram_75__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1771) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5132 ( .A(
        mem_stage_inst_dmem_ram_75__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1772) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5131 ( .A(
        mem_stage_inst_dmem_ram_75__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1773) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5130 ( .A(
        mem_stage_inst_dmem_ram_75__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1774) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5129 ( .A(
        mem_stage_inst_dmem_ram_75__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1775) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5128 ( .A(
        mem_stage_inst_dmem_ram_75__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1776) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5127 ( .A(
        mem_stage_inst_dmem_ram_75__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1777) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5126 ( .A(
        mem_stage_inst_dmem_ram_75__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1778) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5125 ( .A(
        mem_stage_inst_dmem_ram_75__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1779) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5124 ( .A(
        mem_stage_inst_dmem_ram_75__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5914), .Y(mem_stage_inst_dmem_n1780) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5123 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5913) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5122 ( .A(
        mem_stage_inst_dmem_ram_76__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1781) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5121 ( .A(
        mem_stage_inst_dmem_ram_76__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1782) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5120 ( .A(
        mem_stage_inst_dmem_ram_76__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1783) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5119 ( .A(
        mem_stage_inst_dmem_ram_76__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1784) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5118 ( .A(
        mem_stage_inst_dmem_ram_76__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1785) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5117 ( .A(
        mem_stage_inst_dmem_ram_76__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1786) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5116 ( .A(
        mem_stage_inst_dmem_ram_76__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1787) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5115 ( .A(
        mem_stage_inst_dmem_ram_76__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1788) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5114 ( .A(
        mem_stage_inst_dmem_ram_76__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1789) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5113 ( .A(
        mem_stage_inst_dmem_ram_76__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1790) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5112 ( .A(
        mem_stage_inst_dmem_ram_76__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1791) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5111 ( .A(
        mem_stage_inst_dmem_ram_76__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1792) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5110 ( .A(
        mem_stage_inst_dmem_ram_76__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1793) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5109 ( .A(
        mem_stage_inst_dmem_ram_76__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1794) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5108 ( .A(
        mem_stage_inst_dmem_ram_76__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1795) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5107 ( .A(
        mem_stage_inst_dmem_ram_76__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5913), .Y(mem_stage_inst_dmem_n1796) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5106 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5912) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5105 ( .A(
        mem_stage_inst_dmem_ram_77__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1797) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5104 ( .A(
        mem_stage_inst_dmem_ram_77__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1798) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5103 ( .A(
        mem_stage_inst_dmem_ram_77__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1799) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5102 ( .A(
        mem_stage_inst_dmem_ram_77__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1800) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5101 ( .A(
        mem_stage_inst_dmem_ram_77__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1801) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5100 ( .A(
        mem_stage_inst_dmem_ram_77__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1802) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5099 ( .A(
        mem_stage_inst_dmem_ram_77__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1803) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5098 ( .A(
        mem_stage_inst_dmem_ram_77__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1804) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5097 ( .A(
        mem_stage_inst_dmem_ram_77__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1805) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5096 ( .A(
        mem_stage_inst_dmem_ram_77__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1806) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5095 ( .A(
        mem_stage_inst_dmem_ram_77__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1807) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5094 ( .A(
        mem_stage_inst_dmem_ram_77__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1808) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5093 ( .A(
        mem_stage_inst_dmem_ram_77__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1809) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5092 ( .A(
        mem_stage_inst_dmem_ram_77__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1810) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5091 ( .A(
        mem_stage_inst_dmem_ram_77__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1811) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5090 ( .A(
        mem_stage_inst_dmem_ram_77__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5912), .Y(mem_stage_inst_dmem_n1812) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5089 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5911) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5088 ( .A(
        mem_stage_inst_dmem_ram_78__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1813) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5087 ( .A(
        mem_stage_inst_dmem_ram_78__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1814) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5086 ( .A(
        mem_stage_inst_dmem_ram_78__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1815) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5085 ( .A(
        mem_stage_inst_dmem_ram_78__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1816) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5084 ( .A(
        mem_stage_inst_dmem_ram_78__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1817) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5083 ( .A(
        mem_stage_inst_dmem_ram_78__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1818) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5082 ( .A(
        mem_stage_inst_dmem_ram_78__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1819) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5081 ( .A(
        mem_stage_inst_dmem_ram_78__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1820) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5080 ( .A(
        mem_stage_inst_dmem_ram_78__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1821) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5079 ( .A(
        mem_stage_inst_dmem_ram_78__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1822) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5078 ( .A(
        mem_stage_inst_dmem_ram_78__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1823) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5077 ( .A(
        mem_stage_inst_dmem_ram_78__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1824) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5076 ( .A(
        mem_stage_inst_dmem_ram_78__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1825) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5075 ( .A(
        mem_stage_inst_dmem_ram_78__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1826) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5074 ( .A(
        mem_stage_inst_dmem_ram_78__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1827) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5073 ( .A(
        mem_stage_inst_dmem_ram_78__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5911), .Y(mem_stage_inst_dmem_n1828) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5072 ( .A(mem_stage_inst_dmem_n5910), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5909) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5071 ( .A(
        mem_stage_inst_dmem_ram_79__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1829) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5070 ( .A(
        mem_stage_inst_dmem_ram_79__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1830) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5069 ( .A(
        mem_stage_inst_dmem_ram_79__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1831) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5068 ( .A(
        mem_stage_inst_dmem_ram_79__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1832) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5067 ( .A(
        mem_stage_inst_dmem_ram_79__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1833) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5066 ( .A(
        mem_stage_inst_dmem_ram_79__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1834) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5065 ( .A(
        mem_stage_inst_dmem_ram_79__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1835) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5064 ( .A(
        mem_stage_inst_dmem_ram_79__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1836) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5063 ( .A(
        mem_stage_inst_dmem_ram_79__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1837) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5062 ( .A(
        mem_stage_inst_dmem_ram_79__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1838) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5061 ( .A(
        mem_stage_inst_dmem_ram_79__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1839) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5060 ( .A(
        mem_stage_inst_dmem_ram_79__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1840) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5059 ( .A(
        mem_stage_inst_dmem_ram_79__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1841) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5058 ( .A(
        mem_stage_inst_dmem_ram_79__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1842) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5057 ( .A(
        mem_stage_inst_dmem_ram_79__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1843) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5056 ( .A(
        mem_stage_inst_dmem_ram_79__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5909), .Y(mem_stage_inst_dmem_n1844) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5055 ( .A(mem_stage_inst_dmem_n5874), 
        .B(mem_stage_inst_dmem_n5768), .Y(mem_stage_inst_dmem_n5893) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5054 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5908) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5053 ( .A(
        mem_stage_inst_dmem_ram_80__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1845) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5052 ( .A(
        mem_stage_inst_dmem_ram_80__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1846) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5051 ( .A(
        mem_stage_inst_dmem_ram_80__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1847) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5050 ( .A(
        mem_stage_inst_dmem_ram_80__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1848) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5049 ( .A(
        mem_stage_inst_dmem_ram_80__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1849) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5048 ( .A(
        mem_stage_inst_dmem_ram_80__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1850) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5047 ( .A(
        mem_stage_inst_dmem_ram_80__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1851) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5046 ( .A(
        mem_stage_inst_dmem_ram_80__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1852) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5045 ( .A(
        mem_stage_inst_dmem_ram_80__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1853) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5044 ( .A(
        mem_stage_inst_dmem_ram_80__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1854) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5043 ( .A(
        mem_stage_inst_dmem_ram_80__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1855) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5042 ( .A(
        mem_stage_inst_dmem_ram_80__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1856) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5041 ( .A(
        mem_stage_inst_dmem_ram_80__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1857) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5040 ( .A(
        mem_stage_inst_dmem_ram_80__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1858) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5039 ( .A(
        mem_stage_inst_dmem_ram_80__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1859) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5038 ( .A(
        mem_stage_inst_dmem_ram_80__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5908), .Y(mem_stage_inst_dmem_n1860) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5037 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5907) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5036 ( .A(
        mem_stage_inst_dmem_ram_81__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1861) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5035 ( .A(
        mem_stage_inst_dmem_ram_81__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1862) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5034 ( .A(
        mem_stage_inst_dmem_ram_81__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1863) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5033 ( .A(
        mem_stage_inst_dmem_ram_81__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1864) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5032 ( .A(
        mem_stage_inst_dmem_ram_81__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1865) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5031 ( .A(
        mem_stage_inst_dmem_ram_81__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1866) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5030 ( .A(
        mem_stage_inst_dmem_ram_81__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1867) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5029 ( .A(
        mem_stage_inst_dmem_ram_81__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1868) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5028 ( .A(
        mem_stage_inst_dmem_ram_81__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1869) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5027 ( .A(
        mem_stage_inst_dmem_ram_81__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1870) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5026 ( .A(
        mem_stage_inst_dmem_ram_81__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1871) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5025 ( .A(
        mem_stage_inst_dmem_ram_81__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1872) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5024 ( .A(
        mem_stage_inst_dmem_ram_81__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1873) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5023 ( .A(
        mem_stage_inst_dmem_ram_81__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1874) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5022 ( .A(
        mem_stage_inst_dmem_ram_81__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1875) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5021 ( .A(
        mem_stage_inst_dmem_ram_81__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5907), .Y(mem_stage_inst_dmem_n1876) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5020 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5906) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5019 ( .A(
        mem_stage_inst_dmem_ram_82__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1877) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5018 ( .A(
        mem_stage_inst_dmem_ram_82__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1878) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5017 ( .A(
        mem_stage_inst_dmem_ram_82__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1879) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5016 ( .A(
        mem_stage_inst_dmem_ram_82__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1880) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5015 ( .A(
        mem_stage_inst_dmem_ram_82__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1881) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5014 ( .A(
        mem_stage_inst_dmem_ram_82__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1882) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5013 ( .A(
        mem_stage_inst_dmem_ram_82__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1883) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5012 ( .A(
        mem_stage_inst_dmem_ram_82__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1884) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5011 ( .A(
        mem_stage_inst_dmem_ram_82__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1885) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5010 ( .A(
        mem_stage_inst_dmem_ram_82__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1886) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5009 ( .A(
        mem_stage_inst_dmem_ram_82__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1887) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5008 ( .A(
        mem_stage_inst_dmem_ram_82__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1888) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5007 ( .A(
        mem_stage_inst_dmem_ram_82__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1889) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5006 ( .A(
        mem_stage_inst_dmem_ram_82__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1890) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5005 ( .A(
        mem_stage_inst_dmem_ram_82__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1891) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5004 ( .A(
        mem_stage_inst_dmem_ram_82__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5906), .Y(mem_stage_inst_dmem_n1892) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u5003 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5905) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5002 ( .A(
        mem_stage_inst_dmem_ram_83__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1893) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5001 ( .A(
        mem_stage_inst_dmem_ram_83__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1894) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u5000 ( .A(
        mem_stage_inst_dmem_ram_83__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1895) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4999 ( .A(
        mem_stage_inst_dmem_ram_83__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1896) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4998 ( .A(
        mem_stage_inst_dmem_ram_83__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1897) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4997 ( .A(
        mem_stage_inst_dmem_ram_83__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1898) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4996 ( .A(
        mem_stage_inst_dmem_ram_83__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1899) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4995 ( .A(
        mem_stage_inst_dmem_ram_83__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1900) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4994 ( .A(
        mem_stage_inst_dmem_ram_83__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1901) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4993 ( .A(
        mem_stage_inst_dmem_ram_83__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1902) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4992 ( .A(
        mem_stage_inst_dmem_ram_83__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1903) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4991 ( .A(
        mem_stage_inst_dmem_ram_83__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1904) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4990 ( .A(
        mem_stage_inst_dmem_ram_83__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1905) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4989 ( .A(
        mem_stage_inst_dmem_ram_83__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1906) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4988 ( .A(
        mem_stage_inst_dmem_ram_83__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1907) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4987 ( .A(
        mem_stage_inst_dmem_ram_83__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5905), .Y(mem_stage_inst_dmem_n1908) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4986 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5904) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4985 ( .A(
        mem_stage_inst_dmem_ram_84__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1909) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4984 ( .A(
        mem_stage_inst_dmem_ram_84__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1910) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4983 ( .A(
        mem_stage_inst_dmem_ram_84__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1911) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4982 ( .A(
        mem_stage_inst_dmem_ram_84__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1912) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4981 ( .A(
        mem_stage_inst_dmem_ram_84__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1913) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4980 ( .A(
        mem_stage_inst_dmem_ram_84__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1914) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4979 ( .A(
        mem_stage_inst_dmem_ram_84__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1915) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4978 ( .A(
        mem_stage_inst_dmem_ram_84__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1916) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4977 ( .A(
        mem_stage_inst_dmem_ram_84__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1917) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4976 ( .A(
        mem_stage_inst_dmem_ram_84__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1918) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4975 ( .A(
        mem_stage_inst_dmem_ram_84__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1919) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4974 ( .A(
        mem_stage_inst_dmem_ram_84__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1920) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4973 ( .A(
        mem_stage_inst_dmem_ram_84__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1921) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4972 ( .A(
        mem_stage_inst_dmem_ram_84__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1922) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4971 ( .A(
        mem_stage_inst_dmem_ram_84__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1923) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4970 ( .A(
        mem_stage_inst_dmem_ram_84__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5904), .Y(mem_stage_inst_dmem_n1924) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4969 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5903) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4968 ( .A(
        mem_stage_inst_dmem_ram_85__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1925) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4967 ( .A(
        mem_stage_inst_dmem_ram_85__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1926) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4966 ( .A(
        mem_stage_inst_dmem_ram_85__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1927) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4965 ( .A(
        mem_stage_inst_dmem_ram_85__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1928) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4964 ( .A(
        mem_stage_inst_dmem_ram_85__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1929) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4963 ( .A(
        mem_stage_inst_dmem_ram_85__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1930) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4962 ( .A(
        mem_stage_inst_dmem_ram_85__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1931) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4961 ( .A(
        mem_stage_inst_dmem_ram_85__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1932) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4960 ( .A(
        mem_stage_inst_dmem_ram_85__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1933) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4959 ( .A(
        mem_stage_inst_dmem_ram_85__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1934) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4958 ( .A(
        mem_stage_inst_dmem_ram_85__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1935) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4957 ( .A(
        mem_stage_inst_dmem_ram_85__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1936) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4956 ( .A(
        mem_stage_inst_dmem_ram_85__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1937) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4955 ( .A(
        mem_stage_inst_dmem_ram_85__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1938) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4954 ( .A(
        mem_stage_inst_dmem_ram_85__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1939) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4953 ( .A(
        mem_stage_inst_dmem_ram_85__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5903), .Y(mem_stage_inst_dmem_n1940) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4952 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5902) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4951 ( .A(
        mem_stage_inst_dmem_ram_86__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1941) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4950 ( .A(
        mem_stage_inst_dmem_ram_86__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1942) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4949 ( .A(
        mem_stage_inst_dmem_ram_86__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1943) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4948 ( .A(
        mem_stage_inst_dmem_ram_86__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1944) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4947 ( .A(
        mem_stage_inst_dmem_ram_86__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1945) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4946 ( .A(
        mem_stage_inst_dmem_ram_86__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1946) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4945 ( .A(
        mem_stage_inst_dmem_ram_86__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1947) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4944 ( .A(
        mem_stage_inst_dmem_ram_86__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1948) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4943 ( .A(
        mem_stage_inst_dmem_ram_86__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1949) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4942 ( .A(
        mem_stage_inst_dmem_ram_86__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1950) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4941 ( .A(
        mem_stage_inst_dmem_ram_86__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1951) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4940 ( .A(
        mem_stage_inst_dmem_ram_86__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1952) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4939 ( .A(
        mem_stage_inst_dmem_ram_86__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1953) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4938 ( .A(
        mem_stage_inst_dmem_ram_86__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1954) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4937 ( .A(
        mem_stage_inst_dmem_ram_86__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1955) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4936 ( .A(
        mem_stage_inst_dmem_ram_86__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5902), .Y(mem_stage_inst_dmem_n1956) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4935 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5901) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4934 ( .A(
        mem_stage_inst_dmem_ram_87__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1957) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4933 ( .A(
        mem_stage_inst_dmem_ram_87__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1958) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4932 ( .A(
        mem_stage_inst_dmem_ram_87__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1959) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4931 ( .A(
        mem_stage_inst_dmem_ram_87__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1960) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4930 ( .A(
        mem_stage_inst_dmem_ram_87__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1961) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4929 ( .A(
        mem_stage_inst_dmem_ram_87__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1962) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4928 ( .A(
        mem_stage_inst_dmem_ram_87__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1963) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4927 ( .A(
        mem_stage_inst_dmem_ram_87__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1964) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4926 ( .A(
        mem_stage_inst_dmem_ram_87__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1965) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4925 ( .A(
        mem_stage_inst_dmem_ram_87__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1966) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4924 ( .A(
        mem_stage_inst_dmem_ram_87__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1967) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4923 ( .A(
        mem_stage_inst_dmem_ram_87__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1968) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4922 ( .A(
        mem_stage_inst_dmem_ram_87__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1969) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4921 ( .A(
        mem_stage_inst_dmem_ram_87__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1970) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4920 ( .A(
        mem_stage_inst_dmem_ram_87__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1971) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4919 ( .A(
        mem_stage_inst_dmem_ram_87__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5901), .Y(mem_stage_inst_dmem_n1972) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4918 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5900) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4917 ( .A(
        mem_stage_inst_dmem_ram_88__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1973) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4916 ( .A(
        mem_stage_inst_dmem_ram_88__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1974) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4915 ( .A(
        mem_stage_inst_dmem_ram_88__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1975) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4914 ( .A(
        mem_stage_inst_dmem_ram_88__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1976) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4913 ( .A(
        mem_stage_inst_dmem_ram_88__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1977) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4912 ( .A(
        mem_stage_inst_dmem_ram_88__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1978) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4911 ( .A(
        mem_stage_inst_dmem_ram_88__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1979) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4910 ( .A(
        mem_stage_inst_dmem_ram_88__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1980) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4909 ( .A(
        mem_stage_inst_dmem_ram_88__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1981) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4908 ( .A(
        mem_stage_inst_dmem_ram_88__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1982) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4907 ( .A(
        mem_stage_inst_dmem_ram_88__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1983) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4906 ( .A(
        mem_stage_inst_dmem_ram_88__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1984) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4905 ( .A(
        mem_stage_inst_dmem_ram_88__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1985) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4904 ( .A(
        mem_stage_inst_dmem_ram_88__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1986) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4903 ( .A(
        mem_stage_inst_dmem_ram_88__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1987) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4902 ( .A(
        mem_stage_inst_dmem_ram_88__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5900), .Y(mem_stage_inst_dmem_n1988) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4901 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5899) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4900 ( .A(
        mem_stage_inst_dmem_ram_89__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1989) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4899 ( .A(
        mem_stage_inst_dmem_ram_89__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1990) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4898 ( .A(
        mem_stage_inst_dmem_ram_89__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1991) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4897 ( .A(
        mem_stage_inst_dmem_ram_89__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1992) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4896 ( .A(
        mem_stage_inst_dmem_ram_89__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1993) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4895 ( .A(
        mem_stage_inst_dmem_ram_89__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1994) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4894 ( .A(
        mem_stage_inst_dmem_ram_89__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1995) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4893 ( .A(
        mem_stage_inst_dmem_ram_89__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1996) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4892 ( .A(
        mem_stage_inst_dmem_ram_89__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1997) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4891 ( .A(
        mem_stage_inst_dmem_ram_89__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1998) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4890 ( .A(
        mem_stage_inst_dmem_ram_89__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n1999) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4889 ( .A(
        mem_stage_inst_dmem_ram_89__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n2000) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4888 ( .A(
        mem_stage_inst_dmem_ram_89__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n2001) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4887 ( .A(
        mem_stage_inst_dmem_ram_89__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n2002) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4886 ( .A(
        mem_stage_inst_dmem_ram_89__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n2003) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4885 ( .A(
        mem_stage_inst_dmem_ram_89__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5899), .Y(mem_stage_inst_dmem_n2004) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4884 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5898) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4883 ( .A(
        mem_stage_inst_dmem_ram_90__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2005) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4882 ( .A(
        mem_stage_inst_dmem_ram_90__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2006) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4881 ( .A(
        mem_stage_inst_dmem_ram_90__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2007) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4880 ( .A(
        mem_stage_inst_dmem_ram_90__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2008) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4879 ( .A(
        mem_stage_inst_dmem_ram_90__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2009) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4878 ( .A(
        mem_stage_inst_dmem_ram_90__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2010) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4877 ( .A(
        mem_stage_inst_dmem_ram_90__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2011) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4876 ( .A(
        mem_stage_inst_dmem_ram_90__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2012) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4875 ( .A(
        mem_stage_inst_dmem_ram_90__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2013) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4874 ( .A(
        mem_stage_inst_dmem_ram_90__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2014) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4873 ( .A(
        mem_stage_inst_dmem_ram_90__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2015) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4872 ( .A(
        mem_stage_inst_dmem_ram_90__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2016) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4871 ( .A(
        mem_stage_inst_dmem_ram_90__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2017) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4870 ( .A(
        mem_stage_inst_dmem_ram_90__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2018) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4869 ( .A(
        mem_stage_inst_dmem_ram_90__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2019) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4868 ( .A(
        mem_stage_inst_dmem_ram_90__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5898), .Y(mem_stage_inst_dmem_n2020) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4867 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5897) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4866 ( .A(
        mem_stage_inst_dmem_ram_91__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2021) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4865 ( .A(
        mem_stage_inst_dmem_ram_91__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2022) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4864 ( .A(
        mem_stage_inst_dmem_ram_91__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2023) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4863 ( .A(
        mem_stage_inst_dmem_ram_91__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2024) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4862 ( .A(
        mem_stage_inst_dmem_ram_91__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2025) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4861 ( .A(
        mem_stage_inst_dmem_ram_91__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2026) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4860 ( .A(
        mem_stage_inst_dmem_ram_91__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2027) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4859 ( .A(
        mem_stage_inst_dmem_ram_91__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2028) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4858 ( .A(
        mem_stage_inst_dmem_ram_91__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2029) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4857 ( .A(
        mem_stage_inst_dmem_ram_91__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2030) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4856 ( .A(
        mem_stage_inst_dmem_ram_91__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2031) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4855 ( .A(
        mem_stage_inst_dmem_ram_91__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2032) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4854 ( .A(
        mem_stage_inst_dmem_ram_91__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2033) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4853 ( .A(
        mem_stage_inst_dmem_ram_91__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2034) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4852 ( .A(
        mem_stage_inst_dmem_ram_91__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2035) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4851 ( .A(
        mem_stage_inst_dmem_ram_91__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5897), .Y(mem_stage_inst_dmem_n2036) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4850 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5896) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4849 ( .A(
        mem_stage_inst_dmem_ram_92__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2037) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4848 ( .A(
        mem_stage_inst_dmem_ram_92__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2038) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4847 ( .A(
        mem_stage_inst_dmem_ram_92__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2039) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4846 ( .A(
        mem_stage_inst_dmem_ram_92__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2040) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4845 ( .A(
        mem_stage_inst_dmem_ram_92__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2041) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4844 ( .A(
        mem_stage_inst_dmem_ram_92__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2042) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4843 ( .A(
        mem_stage_inst_dmem_ram_92__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2043) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4842 ( .A(
        mem_stage_inst_dmem_ram_92__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2044) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4841 ( .A(
        mem_stage_inst_dmem_ram_92__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2045) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4840 ( .A(
        mem_stage_inst_dmem_ram_92__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2046) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4839 ( .A(
        mem_stage_inst_dmem_ram_92__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2047) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4838 ( .A(
        mem_stage_inst_dmem_ram_92__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2048) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4837 ( .A(
        mem_stage_inst_dmem_ram_92__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2049) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4836 ( .A(
        mem_stage_inst_dmem_ram_92__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2050) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4835 ( .A(
        mem_stage_inst_dmem_ram_92__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2051) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4834 ( .A(
        mem_stage_inst_dmem_ram_92__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5896), .Y(mem_stage_inst_dmem_n2052) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4833 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5895) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4832 ( .A(
        mem_stage_inst_dmem_ram_93__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2053) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4831 ( .A(
        mem_stage_inst_dmem_ram_93__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2054) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4830 ( .A(
        mem_stage_inst_dmem_ram_93__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2055) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4829 ( .A(
        mem_stage_inst_dmem_ram_93__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2056) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4828 ( .A(
        mem_stage_inst_dmem_ram_93__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2057) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4827 ( .A(
        mem_stage_inst_dmem_ram_93__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2058) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4826 ( .A(
        mem_stage_inst_dmem_ram_93__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2059) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4825 ( .A(
        mem_stage_inst_dmem_ram_93__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2060) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4824 ( .A(
        mem_stage_inst_dmem_ram_93__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2061) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4823 ( .A(
        mem_stage_inst_dmem_ram_93__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2062) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4822 ( .A(
        mem_stage_inst_dmem_ram_93__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2063) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4821 ( .A(
        mem_stage_inst_dmem_ram_93__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2064) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4820 ( .A(
        mem_stage_inst_dmem_ram_93__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2065) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4819 ( .A(
        mem_stage_inst_dmem_ram_93__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2066) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4818 ( .A(
        mem_stage_inst_dmem_ram_93__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2067) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4817 ( .A(
        mem_stage_inst_dmem_ram_93__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5895), .Y(mem_stage_inst_dmem_n2068) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4816 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5894) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4815 ( .A(
        mem_stage_inst_dmem_ram_94__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2069) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4814 ( .A(
        mem_stage_inst_dmem_ram_94__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2070) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4813 ( .A(
        mem_stage_inst_dmem_ram_94__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2071) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4812 ( .A(
        mem_stage_inst_dmem_ram_94__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2072) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4811 ( .A(
        mem_stage_inst_dmem_ram_94__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2073) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4810 ( .A(
        mem_stage_inst_dmem_ram_94__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2074) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4809 ( .A(
        mem_stage_inst_dmem_ram_94__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2075) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4808 ( .A(
        mem_stage_inst_dmem_ram_94__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2076) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4807 ( .A(
        mem_stage_inst_dmem_ram_94__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2077) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4806 ( .A(
        mem_stage_inst_dmem_ram_94__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2078) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4805 ( .A(
        mem_stage_inst_dmem_ram_94__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2079) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4804 ( .A(
        mem_stage_inst_dmem_ram_94__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2080) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4803 ( .A(
        mem_stage_inst_dmem_ram_94__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2081) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4802 ( .A(
        mem_stage_inst_dmem_ram_94__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2082) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4801 ( .A(
        mem_stage_inst_dmem_ram_94__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2083) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4800 ( .A(
        mem_stage_inst_dmem_ram_94__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5894), .Y(mem_stage_inst_dmem_n2084) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4799 ( .A(mem_stage_inst_dmem_n5893), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5892) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4798 ( .A(
        mem_stage_inst_dmem_ram_95__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2085) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4797 ( .A(
        mem_stage_inst_dmem_ram_95__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2086) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4796 ( .A(
        mem_stage_inst_dmem_ram_95__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2087) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4795 ( .A(
        mem_stage_inst_dmem_ram_95__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2088) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4794 ( .A(
        mem_stage_inst_dmem_ram_95__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2089) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4793 ( .A(
        mem_stage_inst_dmem_ram_95__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2090) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4792 ( .A(
        mem_stage_inst_dmem_ram_95__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2091) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4791 ( .A(
        mem_stage_inst_dmem_ram_95__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2092) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4790 ( .A(
        mem_stage_inst_dmem_ram_95__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2093) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4789 ( .A(
        mem_stage_inst_dmem_ram_95__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2094) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4788 ( .A(
        mem_stage_inst_dmem_ram_95__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2095) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4787 ( .A(
        mem_stage_inst_dmem_ram_95__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2096) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4786 ( .A(
        mem_stage_inst_dmem_ram_95__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2097) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4785 ( .A(
        mem_stage_inst_dmem_ram_95__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2098) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4784 ( .A(
        mem_stage_inst_dmem_ram_95__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2099) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4783 ( .A(
        mem_stage_inst_dmem_ram_95__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5892), .Y(mem_stage_inst_dmem_n2100) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4782 ( .A(mem_stage_inst_dmem_n5874), 
        .B(mem_stage_inst_dmem_n5750), .Y(mem_stage_inst_dmem_n5876) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4781 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5891) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4780 ( .A(
        mem_stage_inst_dmem_ram_96__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2101) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4779 ( .A(
        mem_stage_inst_dmem_ram_96__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2102) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4778 ( .A(
        mem_stage_inst_dmem_ram_96__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2103) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4777 ( .A(
        mem_stage_inst_dmem_ram_96__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2104) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4776 ( .A(
        mem_stage_inst_dmem_ram_96__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2105) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4775 ( .A(
        mem_stage_inst_dmem_ram_96__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2106) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4774 ( .A(
        mem_stage_inst_dmem_ram_96__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2107) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4773 ( .A(
        mem_stage_inst_dmem_ram_96__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2108) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4772 ( .A(
        mem_stage_inst_dmem_ram_96__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2109) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4771 ( .A(
        mem_stage_inst_dmem_ram_96__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2110) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4770 ( .A(
        mem_stage_inst_dmem_ram_96__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2111) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4769 ( .A(
        mem_stage_inst_dmem_ram_96__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2112) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4768 ( .A(
        mem_stage_inst_dmem_ram_96__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2113) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4767 ( .A(
        mem_stage_inst_dmem_ram_96__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2114) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4766 ( .A(
        mem_stage_inst_dmem_ram_96__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2115) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4765 ( .A(
        mem_stage_inst_dmem_ram_96__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5891), .Y(mem_stage_inst_dmem_n2116) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4764 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5890) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4763 ( .A(
        mem_stage_inst_dmem_ram_97__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2117) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4762 ( .A(
        mem_stage_inst_dmem_ram_97__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2118) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4761 ( .A(
        mem_stage_inst_dmem_ram_97__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2119) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4760 ( .A(
        mem_stage_inst_dmem_ram_97__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2120) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4759 ( .A(
        mem_stage_inst_dmem_ram_97__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2121) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4758 ( .A(
        mem_stage_inst_dmem_ram_97__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2122) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4757 ( .A(
        mem_stage_inst_dmem_ram_97__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2123) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4756 ( .A(
        mem_stage_inst_dmem_ram_97__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2124) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4755 ( .A(
        mem_stage_inst_dmem_ram_97__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2125) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4754 ( .A(
        mem_stage_inst_dmem_ram_97__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2126) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4753 ( .A(
        mem_stage_inst_dmem_ram_97__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2127) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4752 ( .A(
        mem_stage_inst_dmem_ram_97__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2128) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4751 ( .A(
        mem_stage_inst_dmem_ram_97__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2129) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4750 ( .A(
        mem_stage_inst_dmem_ram_97__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2130) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4749 ( .A(
        mem_stage_inst_dmem_ram_97__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2131) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4748 ( .A(
        mem_stage_inst_dmem_ram_97__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5890), .Y(mem_stage_inst_dmem_n2132) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4747 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5889) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4746 ( .A(
        mem_stage_inst_dmem_ram_98__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2133) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4745 ( .A(
        mem_stage_inst_dmem_ram_98__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2134) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4744 ( .A(
        mem_stage_inst_dmem_ram_98__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2135) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4743 ( .A(
        mem_stage_inst_dmem_ram_98__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2136) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4742 ( .A(
        mem_stage_inst_dmem_ram_98__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2137) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4741 ( .A(
        mem_stage_inst_dmem_ram_98__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2138) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4740 ( .A(
        mem_stage_inst_dmem_ram_98__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2139) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4739 ( .A(
        mem_stage_inst_dmem_ram_98__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2140) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4738 ( .A(
        mem_stage_inst_dmem_ram_98__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2141) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4737 ( .A(
        mem_stage_inst_dmem_ram_98__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2142) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4736 ( .A(
        mem_stage_inst_dmem_ram_98__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2143) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4735 ( .A(
        mem_stage_inst_dmem_ram_98__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2144) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4734 ( .A(
        mem_stage_inst_dmem_ram_98__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2145) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4733 ( .A(
        mem_stage_inst_dmem_ram_98__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2146) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4732 ( .A(
        mem_stage_inst_dmem_ram_98__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2147) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4731 ( .A(
        mem_stage_inst_dmem_ram_98__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5889), .Y(mem_stage_inst_dmem_n2148) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4730 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5888) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4729 ( .A(
        mem_stage_inst_dmem_ram_99__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2149) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4728 ( .A(
        mem_stage_inst_dmem_ram_99__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2150) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4727 ( .A(
        mem_stage_inst_dmem_ram_99__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2151) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4726 ( .A(
        mem_stage_inst_dmem_ram_99__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2152) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4725 ( .A(
        mem_stage_inst_dmem_ram_99__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2153) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4724 ( .A(
        mem_stage_inst_dmem_ram_99__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2154) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4723 ( .A(
        mem_stage_inst_dmem_ram_99__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2155) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4722 ( .A(
        mem_stage_inst_dmem_ram_99__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2156) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4721 ( .A(
        mem_stage_inst_dmem_ram_99__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2157) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4720 ( .A(
        mem_stage_inst_dmem_ram_99__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2158) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4719 ( .A(
        mem_stage_inst_dmem_ram_99__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2159) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4718 ( .A(
        mem_stage_inst_dmem_ram_99__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2160) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4717 ( .A(
        mem_stage_inst_dmem_ram_99__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2161) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4716 ( .A(
        mem_stage_inst_dmem_ram_99__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2162) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4715 ( .A(
        mem_stage_inst_dmem_ram_99__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2163) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4714 ( .A(
        mem_stage_inst_dmem_ram_99__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5888), .Y(mem_stage_inst_dmem_n2164) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4713 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5887) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4712 ( .A(
        mem_stage_inst_dmem_ram_100__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2165) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4711 ( .A(
        mem_stage_inst_dmem_ram_100__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2166) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4710 ( .A(
        mem_stage_inst_dmem_ram_100__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2167) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4709 ( .A(
        mem_stage_inst_dmem_ram_100__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2168) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4708 ( .A(
        mem_stage_inst_dmem_ram_100__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2169) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4707 ( .A(
        mem_stage_inst_dmem_ram_100__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2170) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4706 ( .A(
        mem_stage_inst_dmem_ram_100__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2171) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4705 ( .A(
        mem_stage_inst_dmem_ram_100__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2172) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4704 ( .A(
        mem_stage_inst_dmem_ram_100__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2173) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4703 ( .A(
        mem_stage_inst_dmem_ram_100__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2174) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4702 ( .A(
        mem_stage_inst_dmem_ram_100__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2175) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4701 ( .A(
        mem_stage_inst_dmem_ram_100__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2176) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4700 ( .A(
        mem_stage_inst_dmem_ram_100__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2177) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4699 ( .A(
        mem_stage_inst_dmem_ram_100__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2178) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4698 ( .A(
        mem_stage_inst_dmem_ram_100__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2179) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4697 ( .A(
        mem_stage_inst_dmem_ram_100__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5887), .Y(mem_stage_inst_dmem_n2180) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4696 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5886) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4695 ( .A(
        mem_stage_inst_dmem_ram_101__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2181) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4694 ( .A(
        mem_stage_inst_dmem_ram_101__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2182) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4693 ( .A(
        mem_stage_inst_dmem_ram_101__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2183) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4692 ( .A(
        mem_stage_inst_dmem_ram_101__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2184) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4691 ( .A(
        mem_stage_inst_dmem_ram_101__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2185) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4690 ( .A(
        mem_stage_inst_dmem_ram_101__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2186) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4689 ( .A(
        mem_stage_inst_dmem_ram_101__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2187) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4688 ( .A(
        mem_stage_inst_dmem_ram_101__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2188) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4687 ( .A(
        mem_stage_inst_dmem_ram_101__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2189) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4686 ( .A(
        mem_stage_inst_dmem_ram_101__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2190) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4685 ( .A(
        mem_stage_inst_dmem_ram_101__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2191) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4684 ( .A(
        mem_stage_inst_dmem_ram_101__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2192) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4683 ( .A(
        mem_stage_inst_dmem_ram_101__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2193) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4682 ( .A(
        mem_stage_inst_dmem_ram_101__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2194) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4681 ( .A(
        mem_stage_inst_dmem_ram_101__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2195) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4680 ( .A(
        mem_stage_inst_dmem_ram_101__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5886), .Y(mem_stage_inst_dmem_n2196) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4679 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5885) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4678 ( .A(
        mem_stage_inst_dmem_ram_102__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2197) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4677 ( .A(
        mem_stage_inst_dmem_ram_102__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2198) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4676 ( .A(
        mem_stage_inst_dmem_ram_102__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2199) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4675 ( .A(
        mem_stage_inst_dmem_ram_102__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2200) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4674 ( .A(
        mem_stage_inst_dmem_ram_102__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2201) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4673 ( .A(
        mem_stage_inst_dmem_ram_102__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2202) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4672 ( .A(
        mem_stage_inst_dmem_ram_102__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2203) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4671 ( .A(
        mem_stage_inst_dmem_ram_102__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2204) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4670 ( .A(
        mem_stage_inst_dmem_ram_102__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2205) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4669 ( .A(
        mem_stage_inst_dmem_ram_102__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2206) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4668 ( .A(
        mem_stage_inst_dmem_ram_102__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2207) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4667 ( .A(
        mem_stage_inst_dmem_ram_102__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2208) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4666 ( .A(
        mem_stage_inst_dmem_ram_102__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2209) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4665 ( .A(
        mem_stage_inst_dmem_ram_102__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2210) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4664 ( .A(
        mem_stage_inst_dmem_ram_102__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2211) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4663 ( .A(
        mem_stage_inst_dmem_ram_102__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5885), .Y(mem_stage_inst_dmem_n2212) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4662 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5884) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4661 ( .A(
        mem_stage_inst_dmem_ram_103__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2213) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4660 ( .A(
        mem_stage_inst_dmem_ram_103__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2214) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4659 ( .A(
        mem_stage_inst_dmem_ram_103__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2215) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4658 ( .A(
        mem_stage_inst_dmem_ram_103__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2216) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4657 ( .A(
        mem_stage_inst_dmem_ram_103__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2217) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4656 ( .A(
        mem_stage_inst_dmem_ram_103__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2218) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4655 ( .A(
        mem_stage_inst_dmem_ram_103__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2219) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4654 ( .A(
        mem_stage_inst_dmem_ram_103__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2220) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4653 ( .A(
        mem_stage_inst_dmem_ram_103__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2221) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4652 ( .A(
        mem_stage_inst_dmem_ram_103__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2222) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4651 ( .A(
        mem_stage_inst_dmem_ram_103__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2223) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4650 ( .A(
        mem_stage_inst_dmem_ram_103__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2224) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4649 ( .A(
        mem_stage_inst_dmem_ram_103__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2225) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4648 ( .A(
        mem_stage_inst_dmem_ram_103__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2226) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4647 ( .A(
        mem_stage_inst_dmem_ram_103__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2227) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4646 ( .A(
        mem_stage_inst_dmem_ram_103__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5884), .Y(mem_stage_inst_dmem_n2228) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4645 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5883) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4644 ( .A(
        mem_stage_inst_dmem_ram_104__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2229) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4643 ( .A(
        mem_stage_inst_dmem_ram_104__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2230) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4642 ( .A(
        mem_stage_inst_dmem_ram_104__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2231) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4641 ( .A(
        mem_stage_inst_dmem_ram_104__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2232) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4640 ( .A(
        mem_stage_inst_dmem_ram_104__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2233) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4639 ( .A(
        mem_stage_inst_dmem_ram_104__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2234) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4638 ( .A(
        mem_stage_inst_dmem_ram_104__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2235) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4637 ( .A(
        mem_stage_inst_dmem_ram_104__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2236) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4636 ( .A(
        mem_stage_inst_dmem_ram_104__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2237) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4635 ( .A(
        mem_stage_inst_dmem_ram_104__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2238) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4634 ( .A(
        mem_stage_inst_dmem_ram_104__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2239) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4633 ( .A(
        mem_stage_inst_dmem_ram_104__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2240) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4632 ( .A(
        mem_stage_inst_dmem_ram_104__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2241) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4631 ( .A(
        mem_stage_inst_dmem_ram_104__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2242) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4630 ( .A(
        mem_stage_inst_dmem_ram_104__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2243) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4629 ( .A(
        mem_stage_inst_dmem_ram_104__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5883), .Y(mem_stage_inst_dmem_n2244) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4628 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5882) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4627 ( .A(
        mem_stage_inst_dmem_ram_105__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2245) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4626 ( .A(
        mem_stage_inst_dmem_ram_105__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2246) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4625 ( .A(
        mem_stage_inst_dmem_ram_105__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2247) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4624 ( .A(
        mem_stage_inst_dmem_ram_105__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2248) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4623 ( .A(
        mem_stage_inst_dmem_ram_105__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2249) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4622 ( .A(
        mem_stage_inst_dmem_ram_105__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2250) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4621 ( .A(
        mem_stage_inst_dmem_ram_105__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2251) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4620 ( .A(
        mem_stage_inst_dmem_ram_105__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2252) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4619 ( .A(
        mem_stage_inst_dmem_ram_105__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2253) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4618 ( .A(
        mem_stage_inst_dmem_ram_105__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2254) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4617 ( .A(
        mem_stage_inst_dmem_ram_105__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2255) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4616 ( .A(
        mem_stage_inst_dmem_ram_105__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2256) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4615 ( .A(
        mem_stage_inst_dmem_ram_105__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2257) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4614 ( .A(
        mem_stage_inst_dmem_ram_105__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2258) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4613 ( .A(
        mem_stage_inst_dmem_ram_105__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2259) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4612 ( .A(
        mem_stage_inst_dmem_ram_105__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5882), .Y(mem_stage_inst_dmem_n2260) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4611 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5881) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4610 ( .A(
        mem_stage_inst_dmem_ram_106__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2261) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4609 ( .A(
        mem_stage_inst_dmem_ram_106__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2262) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4608 ( .A(
        mem_stage_inst_dmem_ram_106__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2263) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4607 ( .A(
        mem_stage_inst_dmem_ram_106__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2264) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4606 ( .A(
        mem_stage_inst_dmem_ram_106__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2265) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4605 ( .A(
        mem_stage_inst_dmem_ram_106__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2266) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4604 ( .A(
        mem_stage_inst_dmem_ram_106__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2267) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4603 ( .A(
        mem_stage_inst_dmem_ram_106__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2268) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4602 ( .A(
        mem_stage_inst_dmem_ram_106__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2269) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4601 ( .A(
        mem_stage_inst_dmem_ram_106__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2270) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4600 ( .A(
        mem_stage_inst_dmem_ram_106__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2271) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4599 ( .A(
        mem_stage_inst_dmem_ram_106__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2272) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4598 ( .A(
        mem_stage_inst_dmem_ram_106__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2273) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4597 ( .A(
        mem_stage_inst_dmem_ram_106__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2274) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4596 ( .A(
        mem_stage_inst_dmem_ram_106__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2275) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4595 ( .A(
        mem_stage_inst_dmem_ram_106__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5881), .Y(mem_stage_inst_dmem_n2276) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4594 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5880) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4593 ( .A(
        mem_stage_inst_dmem_ram_107__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2277) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4592 ( .A(
        mem_stage_inst_dmem_ram_107__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2278) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4591 ( .A(
        mem_stage_inst_dmem_ram_107__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2279) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4590 ( .A(
        mem_stage_inst_dmem_ram_107__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2280) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4589 ( .A(
        mem_stage_inst_dmem_ram_107__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2281) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4588 ( .A(
        mem_stage_inst_dmem_ram_107__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2282) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4587 ( .A(
        mem_stage_inst_dmem_ram_107__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2283) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4586 ( .A(
        mem_stage_inst_dmem_ram_107__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2284) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4585 ( .A(
        mem_stage_inst_dmem_ram_107__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2285) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4584 ( .A(
        mem_stage_inst_dmem_ram_107__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2286) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4583 ( .A(
        mem_stage_inst_dmem_ram_107__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2287) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4582 ( .A(
        mem_stage_inst_dmem_ram_107__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2288) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4581 ( .A(
        mem_stage_inst_dmem_ram_107__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2289) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4580 ( .A(
        mem_stage_inst_dmem_ram_107__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2290) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4579 ( .A(
        mem_stage_inst_dmem_ram_107__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2291) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4578 ( .A(
        mem_stage_inst_dmem_ram_107__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5880), .Y(mem_stage_inst_dmem_n2292) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4577 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5879) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4576 ( .A(
        mem_stage_inst_dmem_ram_108__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2293) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4575 ( .A(
        mem_stage_inst_dmem_ram_108__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2294) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4574 ( .A(
        mem_stage_inst_dmem_ram_108__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2295) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4573 ( .A(
        mem_stage_inst_dmem_ram_108__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2296) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4572 ( .A(
        mem_stage_inst_dmem_ram_108__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2297) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4571 ( .A(
        mem_stage_inst_dmem_ram_108__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2298) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4570 ( .A(
        mem_stage_inst_dmem_ram_108__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2299) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4569 ( .A(
        mem_stage_inst_dmem_ram_108__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2300) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4568 ( .A(
        mem_stage_inst_dmem_ram_108__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2301) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4567 ( .A(
        mem_stage_inst_dmem_ram_108__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2302) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4566 ( .A(
        mem_stage_inst_dmem_ram_108__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2303) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4565 ( .A(
        mem_stage_inst_dmem_ram_108__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2304) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4564 ( .A(
        mem_stage_inst_dmem_ram_108__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2305) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4563 ( .A(
        mem_stage_inst_dmem_ram_108__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2306) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4562 ( .A(
        mem_stage_inst_dmem_ram_108__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2307) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4561 ( .A(
        mem_stage_inst_dmem_ram_108__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5879), .Y(mem_stage_inst_dmem_n2308) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4560 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5878) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4559 ( .A(
        mem_stage_inst_dmem_ram_109__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2309) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4558 ( .A(
        mem_stage_inst_dmem_ram_109__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2310) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4557 ( .A(
        mem_stage_inst_dmem_ram_109__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2311) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4556 ( .A(
        mem_stage_inst_dmem_ram_109__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2312) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4555 ( .A(
        mem_stage_inst_dmem_ram_109__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2313) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4554 ( .A(
        mem_stage_inst_dmem_ram_109__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2314) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4553 ( .A(
        mem_stage_inst_dmem_ram_109__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2315) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4552 ( .A(
        mem_stage_inst_dmem_ram_109__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2316) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4551 ( .A(
        mem_stage_inst_dmem_ram_109__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2317) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4550 ( .A(
        mem_stage_inst_dmem_ram_109__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2318) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4549 ( .A(
        mem_stage_inst_dmem_ram_109__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2319) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4548 ( .A(
        mem_stage_inst_dmem_ram_109__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2320) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4547 ( .A(
        mem_stage_inst_dmem_ram_109__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2321) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4546 ( .A(
        mem_stage_inst_dmem_ram_109__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2322) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4545 ( .A(
        mem_stage_inst_dmem_ram_109__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2323) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4544 ( .A(
        mem_stage_inst_dmem_ram_109__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5878), .Y(mem_stage_inst_dmem_n2324) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4543 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5877) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4542 ( .A(
        mem_stage_inst_dmem_ram_110__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2325) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4541 ( .A(
        mem_stage_inst_dmem_ram_110__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2326) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4540 ( .A(
        mem_stage_inst_dmem_ram_110__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2327) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4539 ( .A(
        mem_stage_inst_dmem_ram_110__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2328) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4538 ( .A(
        mem_stage_inst_dmem_ram_110__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2329) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4537 ( .A(
        mem_stage_inst_dmem_ram_110__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2330) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4536 ( .A(
        mem_stage_inst_dmem_ram_110__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2331) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4535 ( .A(
        mem_stage_inst_dmem_ram_110__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2332) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4534 ( .A(
        mem_stage_inst_dmem_ram_110__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2333) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4533 ( .A(
        mem_stage_inst_dmem_ram_110__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2334) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4532 ( .A(
        mem_stage_inst_dmem_ram_110__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2335) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4531 ( .A(
        mem_stage_inst_dmem_ram_110__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2336) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4530 ( .A(
        mem_stage_inst_dmem_ram_110__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2337) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4529 ( .A(
        mem_stage_inst_dmem_ram_110__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2338) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4528 ( .A(
        mem_stage_inst_dmem_ram_110__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2339) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4527 ( .A(
        mem_stage_inst_dmem_ram_110__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5877), .Y(mem_stage_inst_dmem_n2340) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4526 ( .A(mem_stage_inst_dmem_n5876), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5875) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4525 ( .A(
        mem_stage_inst_dmem_ram_111__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2341) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4524 ( .A(
        mem_stage_inst_dmem_ram_111__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2342) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4523 ( .A(
        mem_stage_inst_dmem_ram_111__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2343) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4522 ( .A(
        mem_stage_inst_dmem_ram_111__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2344) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4521 ( .A(
        mem_stage_inst_dmem_ram_111__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2345) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4520 ( .A(
        mem_stage_inst_dmem_ram_111__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2346) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4519 ( .A(
        mem_stage_inst_dmem_ram_111__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2347) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4518 ( .A(
        mem_stage_inst_dmem_ram_111__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2348) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4517 ( .A(
        mem_stage_inst_dmem_ram_111__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2349) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4516 ( .A(
        mem_stage_inst_dmem_ram_111__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2350) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4515 ( .A(
        mem_stage_inst_dmem_ram_111__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2351) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4514 ( .A(
        mem_stage_inst_dmem_ram_111__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2352) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4513 ( .A(
        mem_stage_inst_dmem_ram_111__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2353) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4512 ( .A(
        mem_stage_inst_dmem_ram_111__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2354) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4511 ( .A(
        mem_stage_inst_dmem_ram_111__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2355) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4510 ( .A(
        mem_stage_inst_dmem_ram_111__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5875), .Y(mem_stage_inst_dmem_n2356) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4509 ( .A(mem_stage_inst_dmem_n5874), 
        .B(mem_stage_inst_dmem_n5732), .Y(mem_stage_inst_dmem_n5858) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4508 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5873) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4507 ( .A(
        mem_stage_inst_dmem_ram_112__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2357) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4506 ( .A(
        mem_stage_inst_dmem_ram_112__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2358) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4505 ( .A(
        mem_stage_inst_dmem_ram_112__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2359) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4504 ( .A(
        mem_stage_inst_dmem_ram_112__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2360) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4503 ( .A(
        mem_stage_inst_dmem_ram_112__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2361) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4502 ( .A(
        mem_stage_inst_dmem_ram_112__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2362) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4501 ( .A(
        mem_stage_inst_dmem_ram_112__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2363) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4500 ( .A(
        mem_stage_inst_dmem_ram_112__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2364) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4499 ( .A(
        mem_stage_inst_dmem_ram_112__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2365) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4498 ( .A(
        mem_stage_inst_dmem_ram_112__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2366) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4497 ( .A(
        mem_stage_inst_dmem_ram_112__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2367) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4496 ( .A(
        mem_stage_inst_dmem_ram_112__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2368) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4495 ( .A(
        mem_stage_inst_dmem_ram_112__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2369) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4494 ( .A(
        mem_stage_inst_dmem_ram_112__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2370) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4493 ( .A(
        mem_stage_inst_dmem_ram_112__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2371) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4492 ( .A(
        mem_stage_inst_dmem_ram_112__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5873), .Y(mem_stage_inst_dmem_n2372) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4491 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5872) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4490 ( .A(
        mem_stage_inst_dmem_ram_113__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2373) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4489 ( .A(
        mem_stage_inst_dmem_ram_113__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2374) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4488 ( .A(
        mem_stage_inst_dmem_ram_113__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2375) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4487 ( .A(
        mem_stage_inst_dmem_ram_113__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2376) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4486 ( .A(
        mem_stage_inst_dmem_ram_113__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2377) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4485 ( .A(
        mem_stage_inst_dmem_ram_113__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2378) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4484 ( .A(
        mem_stage_inst_dmem_ram_113__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2379) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4483 ( .A(
        mem_stage_inst_dmem_ram_113__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2380) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4482 ( .A(
        mem_stage_inst_dmem_ram_113__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2381) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4481 ( .A(
        mem_stage_inst_dmem_ram_113__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2382) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4480 ( .A(
        mem_stage_inst_dmem_ram_113__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2383) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4479 ( .A(
        mem_stage_inst_dmem_ram_113__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2384) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4478 ( .A(
        mem_stage_inst_dmem_ram_113__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2385) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4477 ( .A(
        mem_stage_inst_dmem_ram_113__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2386) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4476 ( .A(
        mem_stage_inst_dmem_ram_113__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2387) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4475 ( .A(
        mem_stage_inst_dmem_ram_113__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5872), .Y(mem_stage_inst_dmem_n2388) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4474 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5871) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4473 ( .A(
        mem_stage_inst_dmem_ram_114__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2389) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4472 ( .A(
        mem_stage_inst_dmem_ram_114__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2390) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4471 ( .A(
        mem_stage_inst_dmem_ram_114__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2391) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4470 ( .A(
        mem_stage_inst_dmem_ram_114__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2392) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4469 ( .A(
        mem_stage_inst_dmem_ram_114__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2393) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4468 ( .A(
        mem_stage_inst_dmem_ram_114__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2394) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4467 ( .A(
        mem_stage_inst_dmem_ram_114__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2395) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4466 ( .A(
        mem_stage_inst_dmem_ram_114__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2396) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4465 ( .A(
        mem_stage_inst_dmem_ram_114__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2397) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4464 ( .A(
        mem_stage_inst_dmem_ram_114__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2398) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4463 ( .A(
        mem_stage_inst_dmem_ram_114__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2399) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4462 ( .A(
        mem_stage_inst_dmem_ram_114__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2400) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4461 ( .A(
        mem_stage_inst_dmem_ram_114__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2401) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4460 ( .A(
        mem_stage_inst_dmem_ram_114__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2402) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4459 ( .A(
        mem_stage_inst_dmem_ram_114__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2403) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4458 ( .A(
        mem_stage_inst_dmem_ram_114__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5871), .Y(mem_stage_inst_dmem_n2404) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4457 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5870) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4456 ( .A(
        mem_stage_inst_dmem_ram_115__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2405) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4455 ( .A(
        mem_stage_inst_dmem_ram_115__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2406) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4454 ( .A(
        mem_stage_inst_dmem_ram_115__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2407) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4453 ( .A(
        mem_stage_inst_dmem_ram_115__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2408) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4452 ( .A(
        mem_stage_inst_dmem_ram_115__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2409) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4451 ( .A(
        mem_stage_inst_dmem_ram_115__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2410) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4450 ( .A(
        mem_stage_inst_dmem_ram_115__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2411) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4449 ( .A(
        mem_stage_inst_dmem_ram_115__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2412) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4448 ( .A(
        mem_stage_inst_dmem_ram_115__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2413) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4447 ( .A(
        mem_stage_inst_dmem_ram_115__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2414) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4446 ( .A(
        mem_stage_inst_dmem_ram_115__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2415) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4445 ( .A(
        mem_stage_inst_dmem_ram_115__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2416) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4444 ( .A(
        mem_stage_inst_dmem_ram_115__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2417) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4443 ( .A(
        mem_stage_inst_dmem_ram_115__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2418) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4442 ( .A(
        mem_stage_inst_dmem_ram_115__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2419) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4441 ( .A(
        mem_stage_inst_dmem_ram_115__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5870), .Y(mem_stage_inst_dmem_n2420) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4440 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5869) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4439 ( .A(
        mem_stage_inst_dmem_ram_116__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2421) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4438 ( .A(
        mem_stage_inst_dmem_ram_116__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2422) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4437 ( .A(
        mem_stage_inst_dmem_ram_116__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2423) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4436 ( .A(
        mem_stage_inst_dmem_ram_116__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2424) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4435 ( .A(
        mem_stage_inst_dmem_ram_116__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2425) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4434 ( .A(
        mem_stage_inst_dmem_ram_116__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2426) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4433 ( .A(
        mem_stage_inst_dmem_ram_116__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2427) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4432 ( .A(
        mem_stage_inst_dmem_ram_116__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2428) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4431 ( .A(
        mem_stage_inst_dmem_ram_116__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2429) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4430 ( .A(
        mem_stage_inst_dmem_ram_116__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2430) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4429 ( .A(
        mem_stage_inst_dmem_ram_116__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2431) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4428 ( .A(
        mem_stage_inst_dmem_ram_116__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2432) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4427 ( .A(
        mem_stage_inst_dmem_ram_116__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2433) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4426 ( .A(
        mem_stage_inst_dmem_ram_116__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2434) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4425 ( .A(
        mem_stage_inst_dmem_ram_116__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2435) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4424 ( .A(
        mem_stage_inst_dmem_ram_116__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5869), .Y(mem_stage_inst_dmem_n2436) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4423 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5868) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4422 ( .A(
        mem_stage_inst_dmem_ram_117__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2437) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4421 ( .A(
        mem_stage_inst_dmem_ram_117__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2438) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4420 ( .A(
        mem_stage_inst_dmem_ram_117__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2439) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4419 ( .A(
        mem_stage_inst_dmem_ram_117__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2440) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4418 ( .A(
        mem_stage_inst_dmem_ram_117__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2441) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4417 ( .A(
        mem_stage_inst_dmem_ram_117__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2442) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4416 ( .A(
        mem_stage_inst_dmem_ram_117__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2443) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4415 ( .A(
        mem_stage_inst_dmem_ram_117__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2444) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4414 ( .A(
        mem_stage_inst_dmem_ram_117__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2445) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4413 ( .A(
        mem_stage_inst_dmem_ram_117__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2446) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4412 ( .A(
        mem_stage_inst_dmem_ram_117__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2447) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4411 ( .A(
        mem_stage_inst_dmem_ram_117__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2448) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4410 ( .A(
        mem_stage_inst_dmem_ram_117__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2449) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4409 ( .A(
        mem_stage_inst_dmem_ram_117__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2450) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4408 ( .A(
        mem_stage_inst_dmem_ram_117__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2451) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4407 ( .A(
        mem_stage_inst_dmem_ram_117__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5868), .Y(mem_stage_inst_dmem_n2452) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4406 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5867) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4405 ( .A(
        mem_stage_inst_dmem_ram_118__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2453) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4404 ( .A(
        mem_stage_inst_dmem_ram_118__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2454) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4403 ( .A(
        mem_stage_inst_dmem_ram_118__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2455) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4402 ( .A(
        mem_stage_inst_dmem_ram_118__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2456) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4401 ( .A(
        mem_stage_inst_dmem_ram_118__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2457) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4400 ( .A(
        mem_stage_inst_dmem_ram_118__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2458) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4399 ( .A(
        mem_stage_inst_dmem_ram_118__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2459) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4398 ( .A(
        mem_stage_inst_dmem_ram_118__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2460) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4397 ( .A(
        mem_stage_inst_dmem_ram_118__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2461) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4396 ( .A(
        mem_stage_inst_dmem_ram_118__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2462) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4395 ( .A(
        mem_stage_inst_dmem_ram_118__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2463) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4394 ( .A(
        mem_stage_inst_dmem_ram_118__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2464) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4393 ( .A(
        mem_stage_inst_dmem_ram_118__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2465) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4392 ( .A(
        mem_stage_inst_dmem_ram_118__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2466) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4391 ( .A(
        mem_stage_inst_dmem_ram_118__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2467) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4390 ( .A(
        mem_stage_inst_dmem_ram_118__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5867), .Y(mem_stage_inst_dmem_n2468) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4389 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5866) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4388 ( .A(
        mem_stage_inst_dmem_ram_119__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2469) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4387 ( .A(
        mem_stage_inst_dmem_ram_119__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2470) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4386 ( .A(
        mem_stage_inst_dmem_ram_119__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2471) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4385 ( .A(
        mem_stage_inst_dmem_ram_119__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2472) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4384 ( .A(
        mem_stage_inst_dmem_ram_119__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2473) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4383 ( .A(
        mem_stage_inst_dmem_ram_119__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2474) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4382 ( .A(
        mem_stage_inst_dmem_ram_119__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2475) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4381 ( .A(
        mem_stage_inst_dmem_ram_119__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2476) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4380 ( .A(
        mem_stage_inst_dmem_ram_119__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2477) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4379 ( .A(
        mem_stage_inst_dmem_ram_119__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2478) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4378 ( .A(
        mem_stage_inst_dmem_ram_119__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2479) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4377 ( .A(
        mem_stage_inst_dmem_ram_119__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2480) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4376 ( .A(
        mem_stage_inst_dmem_ram_119__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2481) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4375 ( .A(
        mem_stage_inst_dmem_ram_119__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2482) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4374 ( .A(
        mem_stage_inst_dmem_ram_119__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2483) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4373 ( .A(
        mem_stage_inst_dmem_ram_119__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5866), .Y(mem_stage_inst_dmem_n2484) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4372 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5865) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4371 ( .A(
        mem_stage_inst_dmem_ram_120__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2485) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4370 ( .A(
        mem_stage_inst_dmem_ram_120__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2486) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4369 ( .A(
        mem_stage_inst_dmem_ram_120__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2487) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4368 ( .A(
        mem_stage_inst_dmem_ram_120__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2488) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4367 ( .A(
        mem_stage_inst_dmem_ram_120__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2489) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4366 ( .A(
        mem_stage_inst_dmem_ram_120__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2490) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4365 ( .A(
        mem_stage_inst_dmem_ram_120__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2491) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4364 ( .A(
        mem_stage_inst_dmem_ram_120__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2492) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4363 ( .A(
        mem_stage_inst_dmem_ram_120__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2493) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4362 ( .A(
        mem_stage_inst_dmem_ram_120__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2494) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4361 ( .A(
        mem_stage_inst_dmem_ram_120__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2495) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4360 ( .A(
        mem_stage_inst_dmem_ram_120__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2496) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4359 ( .A(
        mem_stage_inst_dmem_ram_120__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2497) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4358 ( .A(
        mem_stage_inst_dmem_ram_120__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2498) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4357 ( .A(
        mem_stage_inst_dmem_ram_120__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2499) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4356 ( .A(
        mem_stage_inst_dmem_ram_120__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5865), .Y(mem_stage_inst_dmem_n2500) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4355 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5864) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4354 ( .A(
        mem_stage_inst_dmem_ram_121__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2501) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4353 ( .A(
        mem_stage_inst_dmem_ram_121__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2502) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4352 ( .A(
        mem_stage_inst_dmem_ram_121__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2503) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4351 ( .A(
        mem_stage_inst_dmem_ram_121__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2504) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4350 ( .A(
        mem_stage_inst_dmem_ram_121__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2505) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4349 ( .A(
        mem_stage_inst_dmem_ram_121__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2506) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4348 ( .A(
        mem_stage_inst_dmem_ram_121__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2507) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4347 ( .A(
        mem_stage_inst_dmem_ram_121__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2508) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4346 ( .A(
        mem_stage_inst_dmem_ram_121__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2509) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4345 ( .A(
        mem_stage_inst_dmem_ram_121__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2510) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4344 ( .A(
        mem_stage_inst_dmem_ram_121__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2511) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4343 ( .A(
        mem_stage_inst_dmem_ram_121__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2512) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4342 ( .A(
        mem_stage_inst_dmem_ram_121__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2513) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4341 ( .A(
        mem_stage_inst_dmem_ram_121__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2514) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4340 ( .A(
        mem_stage_inst_dmem_ram_121__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2515) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4339 ( .A(
        mem_stage_inst_dmem_ram_121__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5864), .Y(mem_stage_inst_dmem_n2516) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4338 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5863) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4337 ( .A(
        mem_stage_inst_dmem_ram_122__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2517) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4336 ( .A(
        mem_stage_inst_dmem_ram_122__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2518) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4335 ( .A(
        mem_stage_inst_dmem_ram_122__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2519) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4334 ( .A(
        mem_stage_inst_dmem_ram_122__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2520) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4333 ( .A(
        mem_stage_inst_dmem_ram_122__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2521) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4332 ( .A(
        mem_stage_inst_dmem_ram_122__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2522) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4331 ( .A(
        mem_stage_inst_dmem_ram_122__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2523) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4330 ( .A(
        mem_stage_inst_dmem_ram_122__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2524) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4329 ( .A(
        mem_stage_inst_dmem_ram_122__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2525) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4328 ( .A(
        mem_stage_inst_dmem_ram_122__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2526) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4327 ( .A(
        mem_stage_inst_dmem_ram_122__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2527) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4326 ( .A(
        mem_stage_inst_dmem_ram_122__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2528) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4325 ( .A(
        mem_stage_inst_dmem_ram_122__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2529) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4324 ( .A(
        mem_stage_inst_dmem_ram_122__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2530) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4323 ( .A(
        mem_stage_inst_dmem_ram_122__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2531) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4322 ( .A(
        mem_stage_inst_dmem_ram_122__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5863), .Y(mem_stage_inst_dmem_n2532) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4321 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5862) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4320 ( .A(
        mem_stage_inst_dmem_ram_123__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2533) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4319 ( .A(
        mem_stage_inst_dmem_ram_123__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2534) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4318 ( .A(
        mem_stage_inst_dmem_ram_123__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2535) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4317 ( .A(
        mem_stage_inst_dmem_ram_123__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2536) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4316 ( .A(
        mem_stage_inst_dmem_ram_123__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2537) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4315 ( .A(
        mem_stage_inst_dmem_ram_123__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2538) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4314 ( .A(
        mem_stage_inst_dmem_ram_123__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2539) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4313 ( .A(
        mem_stage_inst_dmem_ram_123__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2540) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4312 ( .A(
        mem_stage_inst_dmem_ram_123__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2541) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4311 ( .A(
        mem_stage_inst_dmem_ram_123__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2542) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4310 ( .A(
        mem_stage_inst_dmem_ram_123__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2543) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4309 ( .A(
        mem_stage_inst_dmem_ram_123__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2544) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4308 ( .A(
        mem_stage_inst_dmem_ram_123__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2545) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4307 ( .A(
        mem_stage_inst_dmem_ram_123__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2546) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4306 ( .A(
        mem_stage_inst_dmem_ram_123__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2547) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4305 ( .A(
        mem_stage_inst_dmem_ram_123__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5862), .Y(mem_stage_inst_dmem_n2548) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4304 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5861) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4303 ( .A(
        mem_stage_inst_dmem_ram_124__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2549) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4302 ( .A(
        mem_stage_inst_dmem_ram_124__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2550) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4301 ( .A(
        mem_stage_inst_dmem_ram_124__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2551) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4300 ( .A(
        mem_stage_inst_dmem_ram_124__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2552) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4299 ( .A(
        mem_stage_inst_dmem_ram_124__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2553) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4298 ( .A(
        mem_stage_inst_dmem_ram_124__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2554) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4297 ( .A(
        mem_stage_inst_dmem_ram_124__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2555) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4296 ( .A(
        mem_stage_inst_dmem_ram_124__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2556) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4295 ( .A(
        mem_stage_inst_dmem_ram_124__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2557) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4294 ( .A(
        mem_stage_inst_dmem_ram_124__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2558) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4293 ( .A(
        mem_stage_inst_dmem_ram_124__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2559) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4292 ( .A(
        mem_stage_inst_dmem_ram_124__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2560) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4291 ( .A(
        mem_stage_inst_dmem_ram_124__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2561) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4290 ( .A(
        mem_stage_inst_dmem_ram_124__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2562) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4289 ( .A(
        mem_stage_inst_dmem_ram_124__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2563) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4288 ( .A(
        mem_stage_inst_dmem_ram_124__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5861), .Y(mem_stage_inst_dmem_n2564) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4287 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5860) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4286 ( .A(
        mem_stage_inst_dmem_ram_125__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2565) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4285 ( .A(
        mem_stage_inst_dmem_ram_125__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2566) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4284 ( .A(
        mem_stage_inst_dmem_ram_125__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2567) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4283 ( .A(
        mem_stage_inst_dmem_ram_125__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2568) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4282 ( .A(
        mem_stage_inst_dmem_ram_125__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2569) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4281 ( .A(
        mem_stage_inst_dmem_ram_125__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2570) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4280 ( .A(
        mem_stage_inst_dmem_ram_125__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2571) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4279 ( .A(
        mem_stage_inst_dmem_ram_125__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2572) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4278 ( .A(
        mem_stage_inst_dmem_ram_125__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2573) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4277 ( .A(
        mem_stage_inst_dmem_ram_125__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2574) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4276 ( .A(
        mem_stage_inst_dmem_ram_125__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2575) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4275 ( .A(
        mem_stage_inst_dmem_ram_125__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2576) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4274 ( .A(
        mem_stage_inst_dmem_ram_125__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2577) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4273 ( .A(
        mem_stage_inst_dmem_ram_125__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2578) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4272 ( .A(
        mem_stage_inst_dmem_ram_125__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2579) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4271 ( .A(
        mem_stage_inst_dmem_ram_125__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5860), .Y(mem_stage_inst_dmem_n2580) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4270 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5859) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4269 ( .A(
        mem_stage_inst_dmem_ram_126__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2581) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4268 ( .A(
        mem_stage_inst_dmem_ram_126__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2582) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4267 ( .A(
        mem_stage_inst_dmem_ram_126__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2583) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4266 ( .A(
        mem_stage_inst_dmem_ram_126__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2584) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4265 ( .A(
        mem_stage_inst_dmem_ram_126__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2585) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4264 ( .A(
        mem_stage_inst_dmem_ram_126__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2586) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4263 ( .A(
        mem_stage_inst_dmem_ram_126__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2587) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4262 ( .A(
        mem_stage_inst_dmem_ram_126__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2588) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4261 ( .A(
        mem_stage_inst_dmem_ram_126__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2589) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4260 ( .A(
        mem_stage_inst_dmem_ram_126__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2590) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4259 ( .A(
        mem_stage_inst_dmem_ram_126__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2591) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4258 ( .A(
        mem_stage_inst_dmem_ram_126__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2592) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4257 ( .A(
        mem_stage_inst_dmem_ram_126__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2593) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4256 ( .A(
        mem_stage_inst_dmem_ram_126__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2594) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4255 ( .A(
        mem_stage_inst_dmem_ram_126__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2595) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4254 ( .A(
        mem_stage_inst_dmem_ram_126__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5859), .Y(mem_stage_inst_dmem_n2596) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4253 ( .A(mem_stage_inst_dmem_n5858), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5857) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4252 ( .A(
        mem_stage_inst_dmem_ram_127__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2597) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4251 ( .A(
        mem_stage_inst_dmem_ram_127__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2598) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4250 ( .A(
        mem_stage_inst_dmem_ram_127__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2599) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4249 ( .A(
        mem_stage_inst_dmem_ram_127__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2600) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4248 ( .A(
        mem_stage_inst_dmem_ram_127__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2601) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4247 ( .A(
        mem_stage_inst_dmem_ram_127__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2602) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4246 ( .A(
        mem_stage_inst_dmem_ram_127__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2603) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4245 ( .A(
        mem_stage_inst_dmem_ram_127__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2604) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4244 ( .A(
        mem_stage_inst_dmem_ram_127__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2605) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4243 ( .A(
        mem_stage_inst_dmem_ram_127__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2606) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4242 ( .A(
        mem_stage_inst_dmem_ram_127__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2607) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4241 ( .A(
        mem_stage_inst_dmem_ram_127__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2608) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4240 ( .A(
        mem_stage_inst_dmem_ram_127__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2609) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4239 ( .A(
        mem_stage_inst_dmem_ram_127__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2610) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4238 ( .A(
        mem_stage_inst_dmem_ram_127__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2611) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4237 ( .A(
        mem_stage_inst_dmem_ram_127__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5857), .Y(mem_stage_inst_dmem_n2612) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4236 ( .A(ex_pipeline_reg_out[29]), 
        .B(ex_pipeline_reg_out[21]), .Y(mem_stage_inst_dmem_n5786) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4235 ( .A(mem_stage_inst_dmem_n5786), 
        .B(mem_stage_inst_dmem_n5856), .Y(mem_stage_inst_dmem_n5804) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4234 ( .A(mem_stage_inst_dmem_n5804), 
        .B(mem_stage_inst_dmem_n5712), .Y(mem_stage_inst_dmem_n5840) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4233 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5855) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4232 ( .A(
        mem_stage_inst_dmem_ram_128__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2613) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4231 ( .A(
        mem_stage_inst_dmem_ram_128__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2614) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4230 ( .A(
        mem_stage_inst_dmem_ram_128__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2615) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4229 ( .A(
        mem_stage_inst_dmem_ram_128__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2616) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4228 ( .A(
        mem_stage_inst_dmem_ram_128__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2617) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4227 ( .A(
        mem_stage_inst_dmem_ram_128__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2618) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4226 ( .A(
        mem_stage_inst_dmem_ram_128__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2619) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4225 ( .A(
        mem_stage_inst_dmem_ram_128__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2620) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4224 ( .A(
        mem_stage_inst_dmem_ram_128__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2621) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4223 ( .A(
        mem_stage_inst_dmem_ram_128__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2622) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4222 ( .A(
        mem_stage_inst_dmem_ram_128__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2623) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4221 ( .A(
        mem_stage_inst_dmem_ram_128__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2624) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4220 ( .A(
        mem_stage_inst_dmem_ram_128__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2625) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4219 ( .A(
        mem_stage_inst_dmem_ram_128__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2626) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4218 ( .A(
        mem_stage_inst_dmem_ram_128__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2627) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4217 ( .A(
        mem_stage_inst_dmem_ram_128__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5855), .Y(mem_stage_inst_dmem_n2628) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4216 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5854) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4215 ( .A(
        mem_stage_inst_dmem_ram_129__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2629) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4214 ( .A(
        mem_stage_inst_dmem_ram_129__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2630) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4213 ( .A(
        mem_stage_inst_dmem_ram_129__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2631) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4212 ( .A(
        mem_stage_inst_dmem_ram_129__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2632) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4211 ( .A(
        mem_stage_inst_dmem_ram_129__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2633) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4210 ( .A(
        mem_stage_inst_dmem_ram_129__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2634) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4209 ( .A(
        mem_stage_inst_dmem_ram_129__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2635) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4208 ( .A(
        mem_stage_inst_dmem_ram_129__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2636) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4207 ( .A(
        mem_stage_inst_dmem_ram_129__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2637) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4206 ( .A(
        mem_stage_inst_dmem_ram_129__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2638) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4205 ( .A(
        mem_stage_inst_dmem_ram_129__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2639) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4204 ( .A(
        mem_stage_inst_dmem_ram_129__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2640) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4203 ( .A(
        mem_stage_inst_dmem_ram_129__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2641) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4202 ( .A(
        mem_stage_inst_dmem_ram_129__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2642) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4201 ( .A(
        mem_stage_inst_dmem_ram_129__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2643) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4200 ( .A(
        mem_stage_inst_dmem_ram_129__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5854), .Y(mem_stage_inst_dmem_n2644) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4199 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5853) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4198 ( .A(
        mem_stage_inst_dmem_ram_130__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2645) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4197 ( .A(
        mem_stage_inst_dmem_ram_130__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2646) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4196 ( .A(
        mem_stage_inst_dmem_ram_130__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2647) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4195 ( .A(
        mem_stage_inst_dmem_ram_130__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2648) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4194 ( .A(
        mem_stage_inst_dmem_ram_130__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2649) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4193 ( .A(
        mem_stage_inst_dmem_ram_130__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2650) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4192 ( .A(
        mem_stage_inst_dmem_ram_130__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2651) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4191 ( .A(
        mem_stage_inst_dmem_ram_130__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2652) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4190 ( .A(
        mem_stage_inst_dmem_ram_130__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2653) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4189 ( .A(
        mem_stage_inst_dmem_ram_130__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2654) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4188 ( .A(
        mem_stage_inst_dmem_ram_130__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2655) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4187 ( .A(
        mem_stage_inst_dmem_ram_130__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2656) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4186 ( .A(
        mem_stage_inst_dmem_ram_130__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2657) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4185 ( .A(
        mem_stage_inst_dmem_ram_130__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2658) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4184 ( .A(
        mem_stage_inst_dmem_ram_130__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2659) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4183 ( .A(
        mem_stage_inst_dmem_ram_130__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5853), .Y(mem_stage_inst_dmem_n2660) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4182 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5852) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4181 ( .A(
        mem_stage_inst_dmem_ram_131__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2661) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4180 ( .A(
        mem_stage_inst_dmem_ram_131__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2662) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4179 ( .A(
        mem_stage_inst_dmem_ram_131__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2663) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4178 ( .A(
        mem_stage_inst_dmem_ram_131__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2664) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4177 ( .A(
        mem_stage_inst_dmem_ram_131__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2665) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4176 ( .A(
        mem_stage_inst_dmem_ram_131__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2666) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4175 ( .A(
        mem_stage_inst_dmem_ram_131__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2667) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4174 ( .A(
        mem_stage_inst_dmem_ram_131__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2668) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4173 ( .A(
        mem_stage_inst_dmem_ram_131__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2669) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4172 ( .A(
        mem_stage_inst_dmem_ram_131__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2670) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4171 ( .A(
        mem_stage_inst_dmem_ram_131__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2671) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4170 ( .A(
        mem_stage_inst_dmem_ram_131__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2672) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4169 ( .A(
        mem_stage_inst_dmem_ram_131__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2673) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4168 ( .A(
        mem_stage_inst_dmem_ram_131__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2674) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4167 ( .A(
        mem_stage_inst_dmem_ram_131__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2675) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4166 ( .A(
        mem_stage_inst_dmem_ram_131__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5852), .Y(mem_stage_inst_dmem_n2676) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4165 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5851) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4164 ( .A(
        mem_stage_inst_dmem_ram_132__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2677) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4163 ( .A(
        mem_stage_inst_dmem_ram_132__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2678) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4162 ( .A(
        mem_stage_inst_dmem_ram_132__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2679) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4161 ( .A(
        mem_stage_inst_dmem_ram_132__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2680) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4160 ( .A(
        mem_stage_inst_dmem_ram_132__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2681) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4159 ( .A(
        mem_stage_inst_dmem_ram_132__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2682) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4158 ( .A(
        mem_stage_inst_dmem_ram_132__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2683) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4157 ( .A(
        mem_stage_inst_dmem_ram_132__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2684) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4156 ( .A(
        mem_stage_inst_dmem_ram_132__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2685) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4155 ( .A(
        mem_stage_inst_dmem_ram_132__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2686) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4154 ( .A(
        mem_stage_inst_dmem_ram_132__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2687) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4153 ( .A(
        mem_stage_inst_dmem_ram_132__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2688) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4152 ( .A(
        mem_stage_inst_dmem_ram_132__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2689) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4151 ( .A(
        mem_stage_inst_dmem_ram_132__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2690) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4150 ( .A(
        mem_stage_inst_dmem_ram_132__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2691) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4149 ( .A(
        mem_stage_inst_dmem_ram_132__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5851), .Y(mem_stage_inst_dmem_n2692) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4148 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5850) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4147 ( .A(
        mem_stage_inst_dmem_ram_133__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2693) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4146 ( .A(
        mem_stage_inst_dmem_ram_133__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2694) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4145 ( .A(
        mem_stage_inst_dmem_ram_133__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2695) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4144 ( .A(
        mem_stage_inst_dmem_ram_133__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2696) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4143 ( .A(
        mem_stage_inst_dmem_ram_133__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2697) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4142 ( .A(
        mem_stage_inst_dmem_ram_133__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2698) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4141 ( .A(
        mem_stage_inst_dmem_ram_133__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2699) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4140 ( .A(
        mem_stage_inst_dmem_ram_133__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2700) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4139 ( .A(
        mem_stage_inst_dmem_ram_133__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2701) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4138 ( .A(
        mem_stage_inst_dmem_ram_133__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2702) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4137 ( .A(
        mem_stage_inst_dmem_ram_133__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2703) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4136 ( .A(
        mem_stage_inst_dmem_ram_133__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2704) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4135 ( .A(
        mem_stage_inst_dmem_ram_133__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2705) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4134 ( .A(
        mem_stage_inst_dmem_ram_133__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2706) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4133 ( .A(
        mem_stage_inst_dmem_ram_133__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2707) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4132 ( .A(
        mem_stage_inst_dmem_ram_133__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5850), .Y(mem_stage_inst_dmem_n2708) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4131 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5849) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4130 ( .A(
        mem_stage_inst_dmem_ram_134__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2709) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4129 ( .A(
        mem_stage_inst_dmem_ram_134__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2710) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4128 ( .A(
        mem_stage_inst_dmem_ram_134__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2711) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4127 ( .A(
        mem_stage_inst_dmem_ram_134__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2712) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4126 ( .A(
        mem_stage_inst_dmem_ram_134__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2713) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4125 ( .A(
        mem_stage_inst_dmem_ram_134__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2714) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4124 ( .A(
        mem_stage_inst_dmem_ram_134__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2715) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4123 ( .A(
        mem_stage_inst_dmem_ram_134__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2716) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4122 ( .A(
        mem_stage_inst_dmem_ram_134__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2717) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4121 ( .A(
        mem_stage_inst_dmem_ram_134__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2718) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4120 ( .A(
        mem_stage_inst_dmem_ram_134__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2719) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4119 ( .A(
        mem_stage_inst_dmem_ram_134__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2720) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4118 ( .A(
        mem_stage_inst_dmem_ram_134__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2721) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4117 ( .A(
        mem_stage_inst_dmem_ram_134__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2722) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4116 ( .A(
        mem_stage_inst_dmem_ram_134__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2723) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4115 ( .A(
        mem_stage_inst_dmem_ram_134__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5849), .Y(mem_stage_inst_dmem_n2724) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4114 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5848) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4113 ( .A(
        mem_stage_inst_dmem_ram_135__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2725) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4112 ( .A(
        mem_stage_inst_dmem_ram_135__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2726) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4111 ( .A(
        mem_stage_inst_dmem_ram_135__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2727) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4110 ( .A(
        mem_stage_inst_dmem_ram_135__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2728) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4109 ( .A(
        mem_stage_inst_dmem_ram_135__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2729) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4108 ( .A(
        mem_stage_inst_dmem_ram_135__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2730) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4107 ( .A(
        mem_stage_inst_dmem_ram_135__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2731) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4106 ( .A(
        mem_stage_inst_dmem_ram_135__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2732) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4105 ( .A(
        mem_stage_inst_dmem_ram_135__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2733) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4104 ( .A(
        mem_stage_inst_dmem_ram_135__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2734) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4103 ( .A(
        mem_stage_inst_dmem_ram_135__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2735) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4102 ( .A(
        mem_stage_inst_dmem_ram_135__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2736) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4101 ( .A(
        mem_stage_inst_dmem_ram_135__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2737) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4100 ( .A(
        mem_stage_inst_dmem_ram_135__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2738) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4099 ( .A(
        mem_stage_inst_dmem_ram_135__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2739) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4098 ( .A(
        mem_stage_inst_dmem_ram_135__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5848), .Y(mem_stage_inst_dmem_n2740) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4097 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5847) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4096 ( .A(
        mem_stage_inst_dmem_ram_136__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2741) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4095 ( .A(
        mem_stage_inst_dmem_ram_136__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2742) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4094 ( .A(
        mem_stage_inst_dmem_ram_136__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2743) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4093 ( .A(
        mem_stage_inst_dmem_ram_136__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2744) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4092 ( .A(
        mem_stage_inst_dmem_ram_136__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2745) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4091 ( .A(
        mem_stage_inst_dmem_ram_136__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2746) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4090 ( .A(
        mem_stage_inst_dmem_ram_136__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2747) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4089 ( .A(
        mem_stage_inst_dmem_ram_136__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2748) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4088 ( .A(
        mem_stage_inst_dmem_ram_136__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2749) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4087 ( .A(
        mem_stage_inst_dmem_ram_136__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2750) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4086 ( .A(
        mem_stage_inst_dmem_ram_136__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2751) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4085 ( .A(
        mem_stage_inst_dmem_ram_136__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2752) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4084 ( .A(
        mem_stage_inst_dmem_ram_136__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2753) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4083 ( .A(
        mem_stage_inst_dmem_ram_136__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2754) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4082 ( .A(
        mem_stage_inst_dmem_ram_136__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2755) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4081 ( .A(
        mem_stage_inst_dmem_ram_136__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5847), .Y(mem_stage_inst_dmem_n2756) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4080 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5846) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4079 ( .A(
        mem_stage_inst_dmem_ram_137__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2757) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4078 ( .A(
        mem_stage_inst_dmem_ram_137__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2758) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4077 ( .A(
        mem_stage_inst_dmem_ram_137__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2759) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4076 ( .A(
        mem_stage_inst_dmem_ram_137__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2760) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4075 ( .A(
        mem_stage_inst_dmem_ram_137__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2761) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4074 ( .A(
        mem_stage_inst_dmem_ram_137__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2762) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4073 ( .A(
        mem_stage_inst_dmem_ram_137__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2763) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4072 ( .A(
        mem_stage_inst_dmem_ram_137__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2764) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4071 ( .A(
        mem_stage_inst_dmem_ram_137__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2765) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4070 ( .A(
        mem_stage_inst_dmem_ram_137__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2766) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4069 ( .A(
        mem_stage_inst_dmem_ram_137__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2767) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4068 ( .A(
        mem_stage_inst_dmem_ram_137__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2768) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4067 ( .A(
        mem_stage_inst_dmem_ram_137__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2769) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4066 ( .A(
        mem_stage_inst_dmem_ram_137__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2770) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4065 ( .A(
        mem_stage_inst_dmem_ram_137__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2771) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4064 ( .A(
        mem_stage_inst_dmem_ram_137__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5846), .Y(mem_stage_inst_dmem_n2772) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4063 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5845) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4062 ( .A(
        mem_stage_inst_dmem_ram_138__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2773) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4061 ( .A(
        mem_stage_inst_dmem_ram_138__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2774) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4060 ( .A(
        mem_stage_inst_dmem_ram_138__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2775) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4059 ( .A(
        mem_stage_inst_dmem_ram_138__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2776) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4058 ( .A(
        mem_stage_inst_dmem_ram_138__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2777) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4057 ( .A(
        mem_stage_inst_dmem_ram_138__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2778) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4056 ( .A(
        mem_stage_inst_dmem_ram_138__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2779) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4055 ( .A(
        mem_stage_inst_dmem_ram_138__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2780) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4054 ( .A(
        mem_stage_inst_dmem_ram_138__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2781) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4053 ( .A(
        mem_stage_inst_dmem_ram_138__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2782) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4052 ( .A(
        mem_stage_inst_dmem_ram_138__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2783) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4051 ( .A(
        mem_stage_inst_dmem_ram_138__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2784) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4050 ( .A(
        mem_stage_inst_dmem_ram_138__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2785) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4049 ( .A(
        mem_stage_inst_dmem_ram_138__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2786) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4048 ( .A(
        mem_stage_inst_dmem_ram_138__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2787) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4047 ( .A(
        mem_stage_inst_dmem_ram_138__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5845), .Y(mem_stage_inst_dmem_n2788) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4046 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5844) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4045 ( .A(
        mem_stage_inst_dmem_ram_139__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2789) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4044 ( .A(
        mem_stage_inst_dmem_ram_139__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2790) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4043 ( .A(
        mem_stage_inst_dmem_ram_139__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2791) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4042 ( .A(
        mem_stage_inst_dmem_ram_139__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2792) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4041 ( .A(
        mem_stage_inst_dmem_ram_139__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2793) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4040 ( .A(
        mem_stage_inst_dmem_ram_139__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2794) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4039 ( .A(
        mem_stage_inst_dmem_ram_139__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2795) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4038 ( .A(
        mem_stage_inst_dmem_ram_139__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2796) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4037 ( .A(
        mem_stage_inst_dmem_ram_139__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2797) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4036 ( .A(
        mem_stage_inst_dmem_ram_139__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2798) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4035 ( .A(
        mem_stage_inst_dmem_ram_139__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2799) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4034 ( .A(
        mem_stage_inst_dmem_ram_139__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2800) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4033 ( .A(
        mem_stage_inst_dmem_ram_139__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2801) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4032 ( .A(
        mem_stage_inst_dmem_ram_139__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2802) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4031 ( .A(
        mem_stage_inst_dmem_ram_139__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2803) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4030 ( .A(
        mem_stage_inst_dmem_ram_139__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5844), .Y(mem_stage_inst_dmem_n2804) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4029 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5843) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4028 ( .A(
        mem_stage_inst_dmem_ram_140__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2805) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4027 ( .A(
        mem_stage_inst_dmem_ram_140__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2806) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4026 ( .A(
        mem_stage_inst_dmem_ram_140__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2807) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4025 ( .A(
        mem_stage_inst_dmem_ram_140__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2808) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4024 ( .A(
        mem_stage_inst_dmem_ram_140__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2809) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4023 ( .A(
        mem_stage_inst_dmem_ram_140__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2810) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4022 ( .A(
        mem_stage_inst_dmem_ram_140__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2811) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4021 ( .A(
        mem_stage_inst_dmem_ram_140__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2812) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4020 ( .A(
        mem_stage_inst_dmem_ram_140__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2813) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4019 ( .A(
        mem_stage_inst_dmem_ram_140__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2814) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4018 ( .A(
        mem_stage_inst_dmem_ram_140__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2815) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4017 ( .A(
        mem_stage_inst_dmem_ram_140__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2816) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4016 ( .A(
        mem_stage_inst_dmem_ram_140__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2817) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4015 ( .A(
        mem_stage_inst_dmem_ram_140__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2818) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4014 ( .A(
        mem_stage_inst_dmem_ram_140__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2819) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4013 ( .A(
        mem_stage_inst_dmem_ram_140__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5843), .Y(mem_stage_inst_dmem_n2820) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u4012 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5842) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4011 ( .A(
        mem_stage_inst_dmem_ram_141__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2821) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4010 ( .A(
        mem_stage_inst_dmem_ram_141__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2822) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4009 ( .A(
        mem_stage_inst_dmem_ram_141__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2823) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4008 ( .A(
        mem_stage_inst_dmem_ram_141__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2824) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4007 ( .A(
        mem_stage_inst_dmem_ram_141__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2825) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4006 ( .A(
        mem_stage_inst_dmem_ram_141__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2826) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4005 ( .A(
        mem_stage_inst_dmem_ram_141__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2827) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4004 ( .A(
        mem_stage_inst_dmem_ram_141__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2828) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4003 ( .A(
        mem_stage_inst_dmem_ram_141__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2829) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4002 ( .A(
        mem_stage_inst_dmem_ram_141__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2830) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4001 ( .A(
        mem_stage_inst_dmem_ram_141__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2831) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u4000 ( .A(
        mem_stage_inst_dmem_ram_141__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2832) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3999 ( .A(
        mem_stage_inst_dmem_ram_141__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2833) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3998 ( .A(
        mem_stage_inst_dmem_ram_141__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2834) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3997 ( .A(
        mem_stage_inst_dmem_ram_141__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2835) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3996 ( .A(
        mem_stage_inst_dmem_ram_141__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5842), .Y(mem_stage_inst_dmem_n2836) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3995 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5841) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3994 ( .A(
        mem_stage_inst_dmem_ram_142__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2837) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3993 ( .A(
        mem_stage_inst_dmem_ram_142__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2838) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3992 ( .A(
        mem_stage_inst_dmem_ram_142__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2839) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3991 ( .A(
        mem_stage_inst_dmem_ram_142__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2840) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3990 ( .A(
        mem_stage_inst_dmem_ram_142__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2841) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3989 ( .A(
        mem_stage_inst_dmem_ram_142__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2842) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3988 ( .A(
        mem_stage_inst_dmem_ram_142__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2843) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3987 ( .A(
        mem_stage_inst_dmem_ram_142__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2844) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3986 ( .A(
        mem_stage_inst_dmem_ram_142__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2845) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3985 ( .A(
        mem_stage_inst_dmem_ram_142__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2846) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3984 ( .A(
        mem_stage_inst_dmem_ram_142__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2847) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3983 ( .A(
        mem_stage_inst_dmem_ram_142__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2848) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3982 ( .A(
        mem_stage_inst_dmem_ram_142__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2849) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3981 ( .A(
        mem_stage_inst_dmem_ram_142__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2850) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3980 ( .A(
        mem_stage_inst_dmem_ram_142__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2851) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3979 ( .A(
        mem_stage_inst_dmem_ram_142__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5841), .Y(mem_stage_inst_dmem_n2852) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3978 ( .A(mem_stage_inst_dmem_n5840), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5839) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3977 ( .A(
        mem_stage_inst_dmem_ram_143__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2853) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3976 ( .A(
        mem_stage_inst_dmem_ram_143__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2854) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3975 ( .A(
        mem_stage_inst_dmem_ram_143__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2855) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3974 ( .A(
        mem_stage_inst_dmem_ram_143__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2856) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3973 ( .A(
        mem_stage_inst_dmem_ram_143__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2857) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3972 ( .A(
        mem_stage_inst_dmem_ram_143__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2858) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3971 ( .A(
        mem_stage_inst_dmem_ram_143__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2859) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3970 ( .A(
        mem_stage_inst_dmem_ram_143__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2860) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3969 ( .A(
        mem_stage_inst_dmem_ram_143__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2861) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3968 ( .A(
        mem_stage_inst_dmem_ram_143__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2862) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3967 ( .A(
        mem_stage_inst_dmem_ram_143__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2863) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3966 ( .A(
        mem_stage_inst_dmem_ram_143__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2864) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3965 ( .A(
        mem_stage_inst_dmem_ram_143__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2865) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3964 ( .A(
        mem_stage_inst_dmem_ram_143__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2866) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3963 ( .A(
        mem_stage_inst_dmem_ram_143__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2867) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3962 ( .A(
        mem_stage_inst_dmem_ram_143__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5839), .Y(mem_stage_inst_dmem_n2868) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3961 ( .A(mem_stage_inst_dmem_n5804), 
        .B(mem_stage_inst_dmem_n5768), .Y(mem_stage_inst_dmem_n5823) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3960 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5838) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3959 ( .A(
        mem_stage_inst_dmem_ram_144__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2869) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3958 ( .A(
        mem_stage_inst_dmem_ram_144__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2870) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3957 ( .A(
        mem_stage_inst_dmem_ram_144__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2871) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3956 ( .A(
        mem_stage_inst_dmem_ram_144__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2872) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3955 ( .A(
        mem_stage_inst_dmem_ram_144__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2873) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3954 ( .A(
        mem_stage_inst_dmem_ram_144__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2874) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3953 ( .A(
        mem_stage_inst_dmem_ram_144__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2875) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3952 ( .A(
        mem_stage_inst_dmem_ram_144__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2876) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3951 ( .A(
        mem_stage_inst_dmem_ram_144__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2877) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3950 ( .A(
        mem_stage_inst_dmem_ram_144__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2878) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3949 ( .A(
        mem_stage_inst_dmem_ram_144__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2879) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3948 ( .A(
        mem_stage_inst_dmem_ram_144__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2880) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3947 ( .A(
        mem_stage_inst_dmem_ram_144__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2881) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3946 ( .A(
        mem_stage_inst_dmem_ram_144__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2882) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3945 ( .A(
        mem_stage_inst_dmem_ram_144__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2883) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3944 ( .A(
        mem_stage_inst_dmem_ram_144__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5838), .Y(mem_stage_inst_dmem_n2884) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3943 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5837) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3942 ( .A(
        mem_stage_inst_dmem_ram_145__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2885) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3941 ( .A(
        mem_stage_inst_dmem_ram_145__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2886) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3940 ( .A(
        mem_stage_inst_dmem_ram_145__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2887) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3939 ( .A(
        mem_stage_inst_dmem_ram_145__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2888) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3938 ( .A(
        mem_stage_inst_dmem_ram_145__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2889) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3937 ( .A(
        mem_stage_inst_dmem_ram_145__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2890) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3936 ( .A(
        mem_stage_inst_dmem_ram_145__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2891) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3935 ( .A(
        mem_stage_inst_dmem_ram_145__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2892) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3934 ( .A(
        mem_stage_inst_dmem_ram_145__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2893) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3933 ( .A(
        mem_stage_inst_dmem_ram_145__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2894) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3932 ( .A(
        mem_stage_inst_dmem_ram_145__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2895) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3931 ( .A(
        mem_stage_inst_dmem_ram_145__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2896) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3930 ( .A(
        mem_stage_inst_dmem_ram_145__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2897) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3929 ( .A(
        mem_stage_inst_dmem_ram_145__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2898) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3928 ( .A(
        mem_stage_inst_dmem_ram_145__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2899) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3927 ( .A(
        mem_stage_inst_dmem_ram_145__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5837), .Y(mem_stage_inst_dmem_n2900) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3926 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5836) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3925 ( .A(
        mem_stage_inst_dmem_ram_146__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2901) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3924 ( .A(
        mem_stage_inst_dmem_ram_146__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2902) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3923 ( .A(
        mem_stage_inst_dmem_ram_146__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2903) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3922 ( .A(
        mem_stage_inst_dmem_ram_146__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2904) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3921 ( .A(
        mem_stage_inst_dmem_ram_146__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2905) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3920 ( .A(
        mem_stage_inst_dmem_ram_146__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2906) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3919 ( .A(
        mem_stage_inst_dmem_ram_146__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2907) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3918 ( .A(
        mem_stage_inst_dmem_ram_146__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2908) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3917 ( .A(
        mem_stage_inst_dmem_ram_146__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2909) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3916 ( .A(
        mem_stage_inst_dmem_ram_146__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2910) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3915 ( .A(
        mem_stage_inst_dmem_ram_146__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2911) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3914 ( .A(
        mem_stage_inst_dmem_ram_146__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2912) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3913 ( .A(
        mem_stage_inst_dmem_ram_146__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2913) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3912 ( .A(
        mem_stage_inst_dmem_ram_146__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2914) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3911 ( .A(
        mem_stage_inst_dmem_ram_146__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2915) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3910 ( .A(
        mem_stage_inst_dmem_ram_146__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5836), .Y(mem_stage_inst_dmem_n2916) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3909 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5835) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3908 ( .A(
        mem_stage_inst_dmem_ram_147__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2917) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3907 ( .A(
        mem_stage_inst_dmem_ram_147__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2918) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3906 ( .A(
        mem_stage_inst_dmem_ram_147__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2919) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3905 ( .A(
        mem_stage_inst_dmem_ram_147__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2920) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3904 ( .A(
        mem_stage_inst_dmem_ram_147__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2921) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3903 ( .A(
        mem_stage_inst_dmem_ram_147__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2922) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3902 ( .A(
        mem_stage_inst_dmem_ram_147__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2923) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3901 ( .A(
        mem_stage_inst_dmem_ram_147__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2924) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3900 ( .A(
        mem_stage_inst_dmem_ram_147__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2925) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3899 ( .A(
        mem_stage_inst_dmem_ram_147__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2926) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3898 ( .A(
        mem_stage_inst_dmem_ram_147__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2927) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3897 ( .A(
        mem_stage_inst_dmem_ram_147__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2928) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3896 ( .A(
        mem_stage_inst_dmem_ram_147__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2929) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3895 ( .A(
        mem_stage_inst_dmem_ram_147__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2930) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3894 ( .A(
        mem_stage_inst_dmem_ram_147__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2931) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3893 ( .A(
        mem_stage_inst_dmem_ram_147__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5835), .Y(mem_stage_inst_dmem_n2932) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3892 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5834) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3891 ( .A(
        mem_stage_inst_dmem_ram_148__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2933) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3890 ( .A(
        mem_stage_inst_dmem_ram_148__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2934) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3889 ( .A(
        mem_stage_inst_dmem_ram_148__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2935) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3888 ( .A(
        mem_stage_inst_dmem_ram_148__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2936) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3887 ( .A(
        mem_stage_inst_dmem_ram_148__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2937) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3886 ( .A(
        mem_stage_inst_dmem_ram_148__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2938) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3885 ( .A(
        mem_stage_inst_dmem_ram_148__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2939) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3884 ( .A(
        mem_stage_inst_dmem_ram_148__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2940) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3883 ( .A(
        mem_stage_inst_dmem_ram_148__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2941) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3882 ( .A(
        mem_stage_inst_dmem_ram_148__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2942) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3881 ( .A(
        mem_stage_inst_dmem_ram_148__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2943) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3880 ( .A(
        mem_stage_inst_dmem_ram_148__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2944) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3879 ( .A(
        mem_stage_inst_dmem_ram_148__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2945) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3878 ( .A(
        mem_stage_inst_dmem_ram_148__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2946) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3877 ( .A(
        mem_stage_inst_dmem_ram_148__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2947) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3876 ( .A(
        mem_stage_inst_dmem_ram_148__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5834), .Y(mem_stage_inst_dmem_n2948) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3875 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5833) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3874 ( .A(
        mem_stage_inst_dmem_ram_149__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2949) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3873 ( .A(
        mem_stage_inst_dmem_ram_149__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2950) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3872 ( .A(
        mem_stage_inst_dmem_ram_149__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2951) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3871 ( .A(
        mem_stage_inst_dmem_ram_149__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2952) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3870 ( .A(
        mem_stage_inst_dmem_ram_149__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2953) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3869 ( .A(
        mem_stage_inst_dmem_ram_149__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2954) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3868 ( .A(
        mem_stage_inst_dmem_ram_149__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2955) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3867 ( .A(
        mem_stage_inst_dmem_ram_149__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2956) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3866 ( .A(
        mem_stage_inst_dmem_ram_149__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2957) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3865 ( .A(
        mem_stage_inst_dmem_ram_149__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2958) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3864 ( .A(
        mem_stage_inst_dmem_ram_149__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2959) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3863 ( .A(
        mem_stage_inst_dmem_ram_149__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2960) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3862 ( .A(
        mem_stage_inst_dmem_ram_149__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2961) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3861 ( .A(
        mem_stage_inst_dmem_ram_149__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2962) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3860 ( .A(
        mem_stage_inst_dmem_ram_149__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2963) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3859 ( .A(
        mem_stage_inst_dmem_ram_149__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5833), .Y(mem_stage_inst_dmem_n2964) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3858 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5832) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3857 ( .A(
        mem_stage_inst_dmem_ram_150__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2965) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3856 ( .A(
        mem_stage_inst_dmem_ram_150__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2966) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3855 ( .A(
        mem_stage_inst_dmem_ram_150__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2967) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3854 ( .A(
        mem_stage_inst_dmem_ram_150__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2968) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3853 ( .A(
        mem_stage_inst_dmem_ram_150__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2969) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3852 ( .A(
        mem_stage_inst_dmem_ram_150__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2970) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3851 ( .A(
        mem_stage_inst_dmem_ram_150__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2971) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3850 ( .A(
        mem_stage_inst_dmem_ram_150__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2972) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3849 ( .A(
        mem_stage_inst_dmem_ram_150__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2973) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3848 ( .A(
        mem_stage_inst_dmem_ram_150__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2974) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3847 ( .A(
        mem_stage_inst_dmem_ram_150__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2975) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3846 ( .A(
        mem_stage_inst_dmem_ram_150__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2976) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3845 ( .A(
        mem_stage_inst_dmem_ram_150__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2977) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3844 ( .A(
        mem_stage_inst_dmem_ram_150__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2978) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3843 ( .A(
        mem_stage_inst_dmem_ram_150__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2979) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3842 ( .A(
        mem_stage_inst_dmem_ram_150__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5832), .Y(mem_stage_inst_dmem_n2980) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3841 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5831) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3840 ( .A(
        mem_stage_inst_dmem_ram_151__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2981) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3839 ( .A(
        mem_stage_inst_dmem_ram_151__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2982) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3838 ( .A(
        mem_stage_inst_dmem_ram_151__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2983) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3837 ( .A(
        mem_stage_inst_dmem_ram_151__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2984) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3836 ( .A(
        mem_stage_inst_dmem_ram_151__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2985) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3835 ( .A(
        mem_stage_inst_dmem_ram_151__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2986) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3834 ( .A(
        mem_stage_inst_dmem_ram_151__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2987) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3833 ( .A(
        mem_stage_inst_dmem_ram_151__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2988) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3832 ( .A(
        mem_stage_inst_dmem_ram_151__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2989) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3831 ( .A(
        mem_stage_inst_dmem_ram_151__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2990) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3830 ( .A(
        mem_stage_inst_dmem_ram_151__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2991) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3829 ( .A(
        mem_stage_inst_dmem_ram_151__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2992) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3828 ( .A(
        mem_stage_inst_dmem_ram_151__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2993) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3827 ( .A(
        mem_stage_inst_dmem_ram_151__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2994) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3826 ( .A(
        mem_stage_inst_dmem_ram_151__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2995) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3825 ( .A(
        mem_stage_inst_dmem_ram_151__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5831), .Y(mem_stage_inst_dmem_n2996) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3824 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5830) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3823 ( .A(
        mem_stage_inst_dmem_ram_152__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n2997) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3822 ( .A(
        mem_stage_inst_dmem_ram_152__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n2998) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3821 ( .A(
        mem_stage_inst_dmem_ram_152__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n2999) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3820 ( .A(
        mem_stage_inst_dmem_ram_152__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3000) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3819 ( .A(
        mem_stage_inst_dmem_ram_152__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3001) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3818 ( .A(
        mem_stage_inst_dmem_ram_152__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3002) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3817 ( .A(
        mem_stage_inst_dmem_ram_152__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3003) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3816 ( .A(
        mem_stage_inst_dmem_ram_152__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3004) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3815 ( .A(
        mem_stage_inst_dmem_ram_152__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3005) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3814 ( .A(
        mem_stage_inst_dmem_ram_152__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3006) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3813 ( .A(
        mem_stage_inst_dmem_ram_152__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3007) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3812 ( .A(
        mem_stage_inst_dmem_ram_152__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3008) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3811 ( .A(
        mem_stage_inst_dmem_ram_152__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3009) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3810 ( .A(
        mem_stage_inst_dmem_ram_152__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3010) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3809 ( .A(
        mem_stage_inst_dmem_ram_152__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3011) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3808 ( .A(
        mem_stage_inst_dmem_ram_152__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5830), .Y(mem_stage_inst_dmem_n3012) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3807 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5829) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3806 ( .A(
        mem_stage_inst_dmem_ram_153__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3013) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3805 ( .A(
        mem_stage_inst_dmem_ram_153__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3014) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3804 ( .A(
        mem_stage_inst_dmem_ram_153__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3015) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3803 ( .A(
        mem_stage_inst_dmem_ram_153__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3016) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3802 ( .A(
        mem_stage_inst_dmem_ram_153__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3017) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3801 ( .A(
        mem_stage_inst_dmem_ram_153__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3018) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3800 ( .A(
        mem_stage_inst_dmem_ram_153__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3019) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3799 ( .A(
        mem_stage_inst_dmem_ram_153__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3020) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3798 ( .A(
        mem_stage_inst_dmem_ram_153__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3021) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3797 ( .A(
        mem_stage_inst_dmem_ram_153__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3022) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3796 ( .A(
        mem_stage_inst_dmem_ram_153__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3023) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3795 ( .A(
        mem_stage_inst_dmem_ram_153__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3024) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3794 ( .A(
        mem_stage_inst_dmem_ram_153__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3025) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3793 ( .A(
        mem_stage_inst_dmem_ram_153__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3026) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3792 ( .A(
        mem_stage_inst_dmem_ram_153__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3027) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3791 ( .A(
        mem_stage_inst_dmem_ram_153__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5829), .Y(mem_stage_inst_dmem_n3028) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3790 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5828) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3789 ( .A(
        mem_stage_inst_dmem_ram_154__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3029) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3788 ( .A(
        mem_stage_inst_dmem_ram_154__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3030) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3787 ( .A(
        mem_stage_inst_dmem_ram_154__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3031) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3786 ( .A(
        mem_stage_inst_dmem_ram_154__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3032) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3785 ( .A(
        mem_stage_inst_dmem_ram_154__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3033) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3784 ( .A(
        mem_stage_inst_dmem_ram_154__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3034) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3783 ( .A(
        mem_stage_inst_dmem_ram_154__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3035) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3782 ( .A(
        mem_stage_inst_dmem_ram_154__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3036) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3781 ( .A(
        mem_stage_inst_dmem_ram_154__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3037) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3780 ( .A(
        mem_stage_inst_dmem_ram_154__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3038) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3779 ( .A(
        mem_stage_inst_dmem_ram_154__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3039) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3778 ( .A(
        mem_stage_inst_dmem_ram_154__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3040) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3777 ( .A(
        mem_stage_inst_dmem_ram_154__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3041) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3776 ( .A(
        mem_stage_inst_dmem_ram_154__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3042) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3775 ( .A(
        mem_stage_inst_dmem_ram_154__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3043) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3774 ( .A(
        mem_stage_inst_dmem_ram_154__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5828), .Y(mem_stage_inst_dmem_n3044) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3773 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5827) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3772 ( .A(
        mem_stage_inst_dmem_ram_155__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3045) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3771 ( .A(
        mem_stage_inst_dmem_ram_155__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3046) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3770 ( .A(
        mem_stage_inst_dmem_ram_155__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3047) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3769 ( .A(
        mem_stage_inst_dmem_ram_155__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3048) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3768 ( .A(
        mem_stage_inst_dmem_ram_155__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3049) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3767 ( .A(
        mem_stage_inst_dmem_ram_155__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3050) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3766 ( .A(
        mem_stage_inst_dmem_ram_155__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3051) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3765 ( .A(
        mem_stage_inst_dmem_ram_155__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3052) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3764 ( .A(
        mem_stage_inst_dmem_ram_155__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3053) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3763 ( .A(
        mem_stage_inst_dmem_ram_155__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3054) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3762 ( .A(
        mem_stage_inst_dmem_ram_155__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3055) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3761 ( .A(
        mem_stage_inst_dmem_ram_155__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3056) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3760 ( .A(
        mem_stage_inst_dmem_ram_155__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3057) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3759 ( .A(
        mem_stage_inst_dmem_ram_155__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3058) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3758 ( .A(
        mem_stage_inst_dmem_ram_155__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3059) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3757 ( .A(
        mem_stage_inst_dmem_ram_155__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5827), .Y(mem_stage_inst_dmem_n3060) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3756 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5826) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3755 ( .A(
        mem_stage_inst_dmem_ram_156__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3061) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3754 ( .A(
        mem_stage_inst_dmem_ram_156__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3062) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3753 ( .A(
        mem_stage_inst_dmem_ram_156__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3063) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3752 ( .A(
        mem_stage_inst_dmem_ram_156__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3064) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3751 ( .A(
        mem_stage_inst_dmem_ram_156__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3065) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3750 ( .A(
        mem_stage_inst_dmem_ram_156__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3066) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3749 ( .A(
        mem_stage_inst_dmem_ram_156__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3067) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3748 ( .A(
        mem_stage_inst_dmem_ram_156__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3068) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3747 ( .A(
        mem_stage_inst_dmem_ram_156__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3069) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3746 ( .A(
        mem_stage_inst_dmem_ram_156__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3070) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3745 ( .A(
        mem_stage_inst_dmem_ram_156__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3071) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3744 ( .A(
        mem_stage_inst_dmem_ram_156__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3072) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3743 ( .A(
        mem_stage_inst_dmem_ram_156__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3073) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3742 ( .A(
        mem_stage_inst_dmem_ram_156__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3074) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3741 ( .A(
        mem_stage_inst_dmem_ram_156__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3075) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3740 ( .A(
        mem_stage_inst_dmem_ram_156__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5826), .Y(mem_stage_inst_dmem_n3076) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3739 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5825) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3738 ( .A(
        mem_stage_inst_dmem_ram_157__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3077) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3737 ( .A(
        mem_stage_inst_dmem_ram_157__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3078) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3736 ( .A(
        mem_stage_inst_dmem_ram_157__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3079) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3735 ( .A(
        mem_stage_inst_dmem_ram_157__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3080) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3734 ( .A(
        mem_stage_inst_dmem_ram_157__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3081) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3733 ( .A(
        mem_stage_inst_dmem_ram_157__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3082) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3732 ( .A(
        mem_stage_inst_dmem_ram_157__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3083) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3731 ( .A(
        mem_stage_inst_dmem_ram_157__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3084) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3730 ( .A(
        mem_stage_inst_dmem_ram_157__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3085) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3729 ( .A(
        mem_stage_inst_dmem_ram_157__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3086) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3728 ( .A(
        mem_stage_inst_dmem_ram_157__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3087) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3727 ( .A(
        mem_stage_inst_dmem_ram_157__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3088) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3726 ( .A(
        mem_stage_inst_dmem_ram_157__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3089) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3725 ( .A(
        mem_stage_inst_dmem_ram_157__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3090) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3724 ( .A(
        mem_stage_inst_dmem_ram_157__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3091) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3723 ( .A(
        mem_stage_inst_dmem_ram_157__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5825), .Y(mem_stage_inst_dmem_n3092) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3722 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5824) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3721 ( .A(
        mem_stage_inst_dmem_ram_158__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3093) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3720 ( .A(
        mem_stage_inst_dmem_ram_158__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3094) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3719 ( .A(
        mem_stage_inst_dmem_ram_158__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3095) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3718 ( .A(
        mem_stage_inst_dmem_ram_158__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3096) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3717 ( .A(
        mem_stage_inst_dmem_ram_158__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3097) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3716 ( .A(
        mem_stage_inst_dmem_ram_158__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3098) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3715 ( .A(
        mem_stage_inst_dmem_ram_158__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3099) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3714 ( .A(
        mem_stage_inst_dmem_ram_158__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3100) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3713 ( .A(
        mem_stage_inst_dmem_ram_158__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3101) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3712 ( .A(
        mem_stage_inst_dmem_ram_158__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3102) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3711 ( .A(
        mem_stage_inst_dmem_ram_158__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3103) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3710 ( .A(
        mem_stage_inst_dmem_ram_158__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3104) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3709 ( .A(
        mem_stage_inst_dmem_ram_158__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3105) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3708 ( .A(
        mem_stage_inst_dmem_ram_158__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3106) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3707 ( .A(
        mem_stage_inst_dmem_ram_158__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3107) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3706 ( .A(
        mem_stage_inst_dmem_ram_158__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5824), .Y(mem_stage_inst_dmem_n3108) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3705 ( .A(mem_stage_inst_dmem_n5823), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5822) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3704 ( .A(
        mem_stage_inst_dmem_ram_159__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3109) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3703 ( .A(
        mem_stage_inst_dmem_ram_159__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3110) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3702 ( .A(
        mem_stage_inst_dmem_ram_159__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3111) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3701 ( .A(
        mem_stage_inst_dmem_ram_159__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3112) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3700 ( .A(
        mem_stage_inst_dmem_ram_159__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3113) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3699 ( .A(
        mem_stage_inst_dmem_ram_159__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3114) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3698 ( .A(
        mem_stage_inst_dmem_ram_159__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3115) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3697 ( .A(
        mem_stage_inst_dmem_ram_159__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3116) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3696 ( .A(
        mem_stage_inst_dmem_ram_159__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3117) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3695 ( .A(
        mem_stage_inst_dmem_ram_159__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3118) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3694 ( .A(
        mem_stage_inst_dmem_ram_159__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3119) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3693 ( .A(
        mem_stage_inst_dmem_ram_159__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3120) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3692 ( .A(
        mem_stage_inst_dmem_ram_159__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3121) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3691 ( .A(
        mem_stage_inst_dmem_ram_159__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3122) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3690 ( .A(
        mem_stage_inst_dmem_ram_159__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3123) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3689 ( .A(
        mem_stage_inst_dmem_ram_159__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5822), .Y(mem_stage_inst_dmem_n3124) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3688 ( .A(mem_stage_inst_dmem_n5804), 
        .B(mem_stage_inst_dmem_n5750), .Y(mem_stage_inst_dmem_n5806) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3687 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5821) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3686 ( .A(
        mem_stage_inst_dmem_ram_160__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3125) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3685 ( .A(
        mem_stage_inst_dmem_ram_160__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3126) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3684 ( .A(
        mem_stage_inst_dmem_ram_160__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3127) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3683 ( .A(
        mem_stage_inst_dmem_ram_160__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3128) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3682 ( .A(
        mem_stage_inst_dmem_ram_160__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3129) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3681 ( .A(
        mem_stage_inst_dmem_ram_160__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3130) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3680 ( .A(
        mem_stage_inst_dmem_ram_160__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3131) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3679 ( .A(
        mem_stage_inst_dmem_ram_160__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3132) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3678 ( .A(
        mem_stage_inst_dmem_ram_160__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3133) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3677 ( .A(
        mem_stage_inst_dmem_ram_160__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3134) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3676 ( .A(
        mem_stage_inst_dmem_ram_160__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3135) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3675 ( .A(
        mem_stage_inst_dmem_ram_160__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3136) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3674 ( .A(
        mem_stage_inst_dmem_ram_160__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3137) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3673 ( .A(
        mem_stage_inst_dmem_ram_160__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3138) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3672 ( .A(
        mem_stage_inst_dmem_ram_160__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3139) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3671 ( .A(
        mem_stage_inst_dmem_ram_160__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5821), .Y(mem_stage_inst_dmem_n3140) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3670 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5820) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3669 ( .A(
        mem_stage_inst_dmem_ram_161__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3141) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3668 ( .A(
        mem_stage_inst_dmem_ram_161__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3142) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3667 ( .A(
        mem_stage_inst_dmem_ram_161__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3143) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3666 ( .A(
        mem_stage_inst_dmem_ram_161__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3144) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3665 ( .A(
        mem_stage_inst_dmem_ram_161__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3145) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3664 ( .A(
        mem_stage_inst_dmem_ram_161__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3146) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3663 ( .A(
        mem_stage_inst_dmem_ram_161__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3147) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3662 ( .A(
        mem_stage_inst_dmem_ram_161__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3148) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3661 ( .A(
        mem_stage_inst_dmem_ram_161__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3149) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3660 ( .A(
        mem_stage_inst_dmem_ram_161__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3150) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3659 ( .A(
        mem_stage_inst_dmem_ram_161__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3151) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3658 ( .A(
        mem_stage_inst_dmem_ram_161__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3152) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3657 ( .A(
        mem_stage_inst_dmem_ram_161__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3153) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3656 ( .A(
        mem_stage_inst_dmem_ram_161__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3154) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3655 ( .A(
        mem_stage_inst_dmem_ram_161__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3155) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3654 ( .A(
        mem_stage_inst_dmem_ram_161__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5820), .Y(mem_stage_inst_dmem_n3156) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3653 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5819) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3652 ( .A(
        mem_stage_inst_dmem_ram_162__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3157) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3651 ( .A(
        mem_stage_inst_dmem_ram_162__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3158) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3650 ( .A(
        mem_stage_inst_dmem_ram_162__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3159) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3649 ( .A(
        mem_stage_inst_dmem_ram_162__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3160) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3648 ( .A(
        mem_stage_inst_dmem_ram_162__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3161) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3647 ( .A(
        mem_stage_inst_dmem_ram_162__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3162) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3646 ( .A(
        mem_stage_inst_dmem_ram_162__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3163) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3645 ( .A(
        mem_stage_inst_dmem_ram_162__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3164) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3644 ( .A(
        mem_stage_inst_dmem_ram_162__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3165) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3643 ( .A(
        mem_stage_inst_dmem_ram_162__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3166) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3642 ( .A(
        mem_stage_inst_dmem_ram_162__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3167) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3641 ( .A(
        mem_stage_inst_dmem_ram_162__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3168) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3640 ( .A(
        mem_stage_inst_dmem_ram_162__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3169) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3639 ( .A(
        mem_stage_inst_dmem_ram_162__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3170) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3638 ( .A(
        mem_stage_inst_dmem_ram_162__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3171) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3637 ( .A(
        mem_stage_inst_dmem_ram_162__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5819), .Y(mem_stage_inst_dmem_n3172) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3636 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5818) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3635 ( .A(
        mem_stage_inst_dmem_ram_163__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3173) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3634 ( .A(
        mem_stage_inst_dmem_ram_163__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3174) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3633 ( .A(
        mem_stage_inst_dmem_ram_163__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3175) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3632 ( .A(
        mem_stage_inst_dmem_ram_163__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3176) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3631 ( .A(
        mem_stage_inst_dmem_ram_163__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3177) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3630 ( .A(
        mem_stage_inst_dmem_ram_163__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3178) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3629 ( .A(
        mem_stage_inst_dmem_ram_163__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3179) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3628 ( .A(
        mem_stage_inst_dmem_ram_163__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3180) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3627 ( .A(
        mem_stage_inst_dmem_ram_163__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3181) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3626 ( .A(
        mem_stage_inst_dmem_ram_163__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3182) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3625 ( .A(
        mem_stage_inst_dmem_ram_163__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3183) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3624 ( .A(
        mem_stage_inst_dmem_ram_163__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3184) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3623 ( .A(
        mem_stage_inst_dmem_ram_163__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3185) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3622 ( .A(
        mem_stage_inst_dmem_ram_163__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3186) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3621 ( .A(
        mem_stage_inst_dmem_ram_163__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3187) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3620 ( .A(
        mem_stage_inst_dmem_ram_163__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5818), .Y(mem_stage_inst_dmem_n3188) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3619 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5817) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3618 ( .A(
        mem_stage_inst_dmem_ram_164__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3189) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3617 ( .A(
        mem_stage_inst_dmem_ram_164__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3190) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3616 ( .A(
        mem_stage_inst_dmem_ram_164__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3191) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3615 ( .A(
        mem_stage_inst_dmem_ram_164__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3192) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3614 ( .A(
        mem_stage_inst_dmem_ram_164__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3193) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3613 ( .A(
        mem_stage_inst_dmem_ram_164__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3194) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3612 ( .A(
        mem_stage_inst_dmem_ram_164__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3195) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3611 ( .A(
        mem_stage_inst_dmem_ram_164__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3196) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3610 ( .A(
        mem_stage_inst_dmem_ram_164__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3197) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3609 ( .A(
        mem_stage_inst_dmem_ram_164__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3198) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3608 ( .A(
        mem_stage_inst_dmem_ram_164__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3199) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3607 ( .A(
        mem_stage_inst_dmem_ram_164__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3200) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3606 ( .A(
        mem_stage_inst_dmem_ram_164__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3201) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3605 ( .A(
        mem_stage_inst_dmem_ram_164__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3202) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3604 ( .A(
        mem_stage_inst_dmem_ram_164__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3203) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3603 ( .A(
        mem_stage_inst_dmem_ram_164__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5817), .Y(mem_stage_inst_dmem_n3204) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3602 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5816) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3601 ( .A(
        mem_stage_inst_dmem_ram_165__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3205) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3600 ( .A(
        mem_stage_inst_dmem_ram_165__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3206) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3599 ( .A(
        mem_stage_inst_dmem_ram_165__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3207) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3598 ( .A(
        mem_stage_inst_dmem_ram_165__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3208) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3597 ( .A(
        mem_stage_inst_dmem_ram_165__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3209) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3596 ( .A(
        mem_stage_inst_dmem_ram_165__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3210) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3595 ( .A(
        mem_stage_inst_dmem_ram_165__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3211) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3594 ( .A(
        mem_stage_inst_dmem_ram_165__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3212) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3593 ( .A(
        mem_stage_inst_dmem_ram_165__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3213) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3592 ( .A(
        mem_stage_inst_dmem_ram_165__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3214) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3591 ( .A(
        mem_stage_inst_dmem_ram_165__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3215) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3590 ( .A(
        mem_stage_inst_dmem_ram_165__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3216) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3589 ( .A(
        mem_stage_inst_dmem_ram_165__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3217) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3588 ( .A(
        mem_stage_inst_dmem_ram_165__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3218) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3587 ( .A(
        mem_stage_inst_dmem_ram_165__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3219) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3586 ( .A(
        mem_stage_inst_dmem_ram_165__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5816), .Y(mem_stage_inst_dmem_n3220) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3585 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5815) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3584 ( .A(
        mem_stage_inst_dmem_ram_166__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3221) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3583 ( .A(
        mem_stage_inst_dmem_ram_166__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3222) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3582 ( .A(
        mem_stage_inst_dmem_ram_166__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3223) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3581 ( .A(
        mem_stage_inst_dmem_ram_166__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3224) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3580 ( .A(
        mem_stage_inst_dmem_ram_166__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3225) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3579 ( .A(
        mem_stage_inst_dmem_ram_166__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3226) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3578 ( .A(
        mem_stage_inst_dmem_ram_166__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3227) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3577 ( .A(
        mem_stage_inst_dmem_ram_166__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3228) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3576 ( .A(
        mem_stage_inst_dmem_ram_166__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3229) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3575 ( .A(
        mem_stage_inst_dmem_ram_166__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3230) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3574 ( .A(
        mem_stage_inst_dmem_ram_166__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3231) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3573 ( .A(
        mem_stage_inst_dmem_ram_166__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3232) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3572 ( .A(
        mem_stage_inst_dmem_ram_166__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3233) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3571 ( .A(
        mem_stage_inst_dmem_ram_166__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3234) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3570 ( .A(
        mem_stage_inst_dmem_ram_166__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3235) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3569 ( .A(
        mem_stage_inst_dmem_ram_166__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5815), .Y(mem_stage_inst_dmem_n3236) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3568 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5814) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3567 ( .A(
        mem_stage_inst_dmem_ram_167__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3237) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3566 ( .A(
        mem_stage_inst_dmem_ram_167__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3238) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3565 ( .A(
        mem_stage_inst_dmem_ram_167__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3239) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3564 ( .A(
        mem_stage_inst_dmem_ram_167__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3240) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3563 ( .A(
        mem_stage_inst_dmem_ram_167__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3241) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3562 ( .A(
        mem_stage_inst_dmem_ram_167__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3242) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3561 ( .A(
        mem_stage_inst_dmem_ram_167__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3243) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3560 ( .A(
        mem_stage_inst_dmem_ram_167__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3244) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3559 ( .A(
        mem_stage_inst_dmem_ram_167__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3245) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3558 ( .A(
        mem_stage_inst_dmem_ram_167__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3246) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3557 ( .A(
        mem_stage_inst_dmem_ram_167__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3247) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3556 ( .A(
        mem_stage_inst_dmem_ram_167__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3248) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3555 ( .A(
        mem_stage_inst_dmem_ram_167__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3249) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3554 ( .A(
        mem_stage_inst_dmem_ram_167__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3250) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3553 ( .A(
        mem_stage_inst_dmem_ram_167__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3251) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3552 ( .A(
        mem_stage_inst_dmem_ram_167__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5814), .Y(mem_stage_inst_dmem_n3252) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3551 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5813) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3550 ( .A(
        mem_stage_inst_dmem_ram_168__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3253) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3549 ( .A(
        mem_stage_inst_dmem_ram_168__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3254) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3548 ( .A(
        mem_stage_inst_dmem_ram_168__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3255) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3547 ( .A(
        mem_stage_inst_dmem_ram_168__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3256) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3546 ( .A(
        mem_stage_inst_dmem_ram_168__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3257) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3545 ( .A(
        mem_stage_inst_dmem_ram_168__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3258) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3544 ( .A(
        mem_stage_inst_dmem_ram_168__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3259) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3543 ( .A(
        mem_stage_inst_dmem_ram_168__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3260) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3542 ( .A(
        mem_stage_inst_dmem_ram_168__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3261) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3541 ( .A(
        mem_stage_inst_dmem_ram_168__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3262) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3540 ( .A(
        mem_stage_inst_dmem_ram_168__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3263) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3539 ( .A(
        mem_stage_inst_dmem_ram_168__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3264) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3538 ( .A(
        mem_stage_inst_dmem_ram_168__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3265) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3537 ( .A(
        mem_stage_inst_dmem_ram_168__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3266) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3536 ( .A(
        mem_stage_inst_dmem_ram_168__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3267) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3535 ( .A(
        mem_stage_inst_dmem_ram_168__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5813), .Y(mem_stage_inst_dmem_n3268) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3534 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5812) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3533 ( .A(
        mem_stage_inst_dmem_ram_169__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3269) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3532 ( .A(
        mem_stage_inst_dmem_ram_169__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3270) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3531 ( .A(
        mem_stage_inst_dmem_ram_169__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3271) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3530 ( .A(
        mem_stage_inst_dmem_ram_169__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3272) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3529 ( .A(
        mem_stage_inst_dmem_ram_169__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3273) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3528 ( .A(
        mem_stage_inst_dmem_ram_169__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3274) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3527 ( .A(
        mem_stage_inst_dmem_ram_169__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3275) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3526 ( .A(
        mem_stage_inst_dmem_ram_169__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3276) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3525 ( .A(
        mem_stage_inst_dmem_ram_169__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3277) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3524 ( .A(
        mem_stage_inst_dmem_ram_169__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3278) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3523 ( .A(
        mem_stage_inst_dmem_ram_169__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3279) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3522 ( .A(
        mem_stage_inst_dmem_ram_169__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3280) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3521 ( .A(
        mem_stage_inst_dmem_ram_169__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3281) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3520 ( .A(
        mem_stage_inst_dmem_ram_169__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3282) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3519 ( .A(
        mem_stage_inst_dmem_ram_169__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3283) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3518 ( .A(
        mem_stage_inst_dmem_ram_169__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5812), .Y(mem_stage_inst_dmem_n3284) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3517 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5811) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3516 ( .A(
        mem_stage_inst_dmem_ram_170__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3285) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3515 ( .A(
        mem_stage_inst_dmem_ram_170__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3286) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3514 ( .A(
        mem_stage_inst_dmem_ram_170__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3287) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3513 ( .A(
        mem_stage_inst_dmem_ram_170__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3288) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3512 ( .A(
        mem_stage_inst_dmem_ram_170__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3289) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3511 ( .A(
        mem_stage_inst_dmem_ram_170__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3290) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3510 ( .A(
        mem_stage_inst_dmem_ram_170__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3291) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3509 ( .A(
        mem_stage_inst_dmem_ram_170__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3292) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3508 ( .A(
        mem_stage_inst_dmem_ram_170__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3293) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3507 ( .A(
        mem_stage_inst_dmem_ram_170__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3294) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3506 ( .A(
        mem_stage_inst_dmem_ram_170__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3295) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3505 ( .A(
        mem_stage_inst_dmem_ram_170__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3296) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3504 ( .A(
        mem_stage_inst_dmem_ram_170__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3297) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3503 ( .A(
        mem_stage_inst_dmem_ram_170__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3298) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3502 ( .A(
        mem_stage_inst_dmem_ram_170__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3299) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3501 ( .A(
        mem_stage_inst_dmem_ram_170__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5811), .Y(mem_stage_inst_dmem_n3300) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3500 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5810) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3499 ( .A(
        mem_stage_inst_dmem_ram_171__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3301) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3498 ( .A(
        mem_stage_inst_dmem_ram_171__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3302) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3497 ( .A(
        mem_stage_inst_dmem_ram_171__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3303) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3496 ( .A(
        mem_stage_inst_dmem_ram_171__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3304) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3495 ( .A(
        mem_stage_inst_dmem_ram_171__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3305) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3494 ( .A(
        mem_stage_inst_dmem_ram_171__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3306) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3493 ( .A(
        mem_stage_inst_dmem_ram_171__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3307) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3492 ( .A(
        mem_stage_inst_dmem_ram_171__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3308) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3491 ( .A(
        mem_stage_inst_dmem_ram_171__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3309) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3490 ( .A(
        mem_stage_inst_dmem_ram_171__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3310) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3489 ( .A(
        mem_stage_inst_dmem_ram_171__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3311) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3488 ( .A(
        mem_stage_inst_dmem_ram_171__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3312) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3487 ( .A(
        mem_stage_inst_dmem_ram_171__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3313) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3486 ( .A(
        mem_stage_inst_dmem_ram_171__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3314) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3485 ( .A(
        mem_stage_inst_dmem_ram_171__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3315) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3484 ( .A(
        mem_stage_inst_dmem_ram_171__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5810), .Y(mem_stage_inst_dmem_n3316) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3483 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5809) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3482 ( .A(
        mem_stage_inst_dmem_ram_172__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3317) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3481 ( .A(
        mem_stage_inst_dmem_ram_172__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3318) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3480 ( .A(
        mem_stage_inst_dmem_ram_172__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3319) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3479 ( .A(
        mem_stage_inst_dmem_ram_172__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3320) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3478 ( .A(
        mem_stage_inst_dmem_ram_172__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3321) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3477 ( .A(
        mem_stage_inst_dmem_ram_172__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3322) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3476 ( .A(
        mem_stage_inst_dmem_ram_172__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3323) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3475 ( .A(
        mem_stage_inst_dmem_ram_172__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3324) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3474 ( .A(
        mem_stage_inst_dmem_ram_172__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3325) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3473 ( .A(
        mem_stage_inst_dmem_ram_172__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3326) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3472 ( .A(
        mem_stage_inst_dmem_ram_172__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3327) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3471 ( .A(
        mem_stage_inst_dmem_ram_172__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3328) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3470 ( .A(
        mem_stage_inst_dmem_ram_172__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3329) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3469 ( .A(
        mem_stage_inst_dmem_ram_172__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3330) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3468 ( .A(
        mem_stage_inst_dmem_ram_172__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3331) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3467 ( .A(
        mem_stage_inst_dmem_ram_172__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5809), .Y(mem_stage_inst_dmem_n3332) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3466 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5808) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3465 ( .A(
        mem_stage_inst_dmem_ram_173__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3333) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3464 ( .A(
        mem_stage_inst_dmem_ram_173__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3334) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3463 ( .A(
        mem_stage_inst_dmem_ram_173__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3335) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3462 ( .A(
        mem_stage_inst_dmem_ram_173__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3336) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3461 ( .A(
        mem_stage_inst_dmem_ram_173__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3337) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3460 ( .A(
        mem_stage_inst_dmem_ram_173__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3338) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3459 ( .A(
        mem_stage_inst_dmem_ram_173__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3339) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3458 ( .A(
        mem_stage_inst_dmem_ram_173__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3340) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3457 ( .A(
        mem_stage_inst_dmem_ram_173__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3341) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3456 ( .A(
        mem_stage_inst_dmem_ram_173__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3342) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3455 ( .A(
        mem_stage_inst_dmem_ram_173__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3343) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3454 ( .A(
        mem_stage_inst_dmem_ram_173__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3344) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3453 ( .A(
        mem_stage_inst_dmem_ram_173__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3345) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3452 ( .A(
        mem_stage_inst_dmem_ram_173__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3346) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3451 ( .A(
        mem_stage_inst_dmem_ram_173__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3347) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3450 ( .A(
        mem_stage_inst_dmem_ram_173__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5808), .Y(mem_stage_inst_dmem_n3348) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3449 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5807) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3448 ( .A(
        mem_stage_inst_dmem_ram_174__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3349) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3447 ( .A(
        mem_stage_inst_dmem_ram_174__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3350) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3446 ( .A(
        mem_stage_inst_dmem_ram_174__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3351) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3445 ( .A(
        mem_stage_inst_dmem_ram_174__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3352) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3444 ( .A(
        mem_stage_inst_dmem_ram_174__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3353) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3443 ( .A(
        mem_stage_inst_dmem_ram_174__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3354) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3442 ( .A(
        mem_stage_inst_dmem_ram_174__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3355) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3441 ( .A(
        mem_stage_inst_dmem_ram_174__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3356) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3440 ( .A(
        mem_stage_inst_dmem_ram_174__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3357) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3439 ( .A(
        mem_stage_inst_dmem_ram_174__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3358) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3438 ( .A(
        mem_stage_inst_dmem_ram_174__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3359) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3437 ( .A(
        mem_stage_inst_dmem_ram_174__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3360) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3436 ( .A(
        mem_stage_inst_dmem_ram_174__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3361) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3435 ( .A(
        mem_stage_inst_dmem_ram_174__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3362) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3434 ( .A(
        mem_stage_inst_dmem_ram_174__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3363) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3433 ( .A(
        mem_stage_inst_dmem_ram_174__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5807), .Y(mem_stage_inst_dmem_n3364) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3432 ( .A(mem_stage_inst_dmem_n5806), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5805) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3431 ( .A(
        mem_stage_inst_dmem_ram_175__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3365) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3430 ( .A(
        mem_stage_inst_dmem_ram_175__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3366) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3429 ( .A(
        mem_stage_inst_dmem_ram_175__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3367) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3428 ( .A(
        mem_stage_inst_dmem_ram_175__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3368) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3427 ( .A(
        mem_stage_inst_dmem_ram_175__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3369) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3426 ( .A(
        mem_stage_inst_dmem_ram_175__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3370) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3425 ( .A(
        mem_stage_inst_dmem_ram_175__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3371) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3424 ( .A(
        mem_stage_inst_dmem_ram_175__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3372) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3423 ( .A(
        mem_stage_inst_dmem_ram_175__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3373) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3422 ( .A(
        mem_stage_inst_dmem_ram_175__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3374) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3421 ( .A(
        mem_stage_inst_dmem_ram_175__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3375) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3420 ( .A(
        mem_stage_inst_dmem_ram_175__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3376) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3419 ( .A(
        mem_stage_inst_dmem_ram_175__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3377) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3418 ( .A(
        mem_stage_inst_dmem_ram_175__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3378) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3417 ( .A(
        mem_stage_inst_dmem_ram_175__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3379) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3416 ( .A(
        mem_stage_inst_dmem_ram_175__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5805), .Y(mem_stage_inst_dmem_n3380) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3415 ( .A(mem_stage_inst_dmem_n5804), 
        .B(mem_stage_inst_dmem_n5732), .Y(mem_stage_inst_dmem_n5788) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3414 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5803) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3413 ( .A(
        mem_stage_inst_dmem_ram_176__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3381) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3412 ( .A(
        mem_stage_inst_dmem_ram_176__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3382) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3411 ( .A(
        mem_stage_inst_dmem_ram_176__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3383) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3410 ( .A(
        mem_stage_inst_dmem_ram_176__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3384) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3409 ( .A(
        mem_stage_inst_dmem_ram_176__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3385) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3408 ( .A(
        mem_stage_inst_dmem_ram_176__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3386) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3407 ( .A(
        mem_stage_inst_dmem_ram_176__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3387) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3406 ( .A(
        mem_stage_inst_dmem_ram_176__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3388) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3405 ( .A(
        mem_stage_inst_dmem_ram_176__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3389) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3404 ( .A(
        mem_stage_inst_dmem_ram_176__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3390) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3403 ( .A(
        mem_stage_inst_dmem_ram_176__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3391) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3402 ( .A(
        mem_stage_inst_dmem_ram_176__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3392) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3401 ( .A(
        mem_stage_inst_dmem_ram_176__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3393) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3400 ( .A(
        mem_stage_inst_dmem_ram_176__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3394) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3399 ( .A(
        mem_stage_inst_dmem_ram_176__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3395) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3398 ( .A(
        mem_stage_inst_dmem_ram_176__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5803), .Y(mem_stage_inst_dmem_n3396) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3397 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5802) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3396 ( .A(
        mem_stage_inst_dmem_ram_177__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3397) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3395 ( .A(
        mem_stage_inst_dmem_ram_177__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3398) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3394 ( .A(
        mem_stage_inst_dmem_ram_177__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3399) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3393 ( .A(
        mem_stage_inst_dmem_ram_177__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3400) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3392 ( .A(
        mem_stage_inst_dmem_ram_177__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3401) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3391 ( .A(
        mem_stage_inst_dmem_ram_177__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3402) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3390 ( .A(
        mem_stage_inst_dmem_ram_177__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3403) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3389 ( .A(
        mem_stage_inst_dmem_ram_177__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3404) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3388 ( .A(
        mem_stage_inst_dmem_ram_177__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3405) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3387 ( .A(
        mem_stage_inst_dmem_ram_177__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3406) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3386 ( .A(
        mem_stage_inst_dmem_ram_177__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3407) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3385 ( .A(
        mem_stage_inst_dmem_ram_177__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3408) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3384 ( .A(
        mem_stage_inst_dmem_ram_177__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3409) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3383 ( .A(
        mem_stage_inst_dmem_ram_177__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3410) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3382 ( .A(
        mem_stage_inst_dmem_ram_177__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3411) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3381 ( .A(
        mem_stage_inst_dmem_ram_177__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5802), .Y(mem_stage_inst_dmem_n3412) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3380 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5801) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3379 ( .A(
        mem_stage_inst_dmem_ram_178__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3413) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3378 ( .A(
        mem_stage_inst_dmem_ram_178__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3414) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3377 ( .A(
        mem_stage_inst_dmem_ram_178__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3415) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3376 ( .A(
        mem_stage_inst_dmem_ram_178__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3416) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3375 ( .A(
        mem_stage_inst_dmem_ram_178__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3417) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3374 ( .A(
        mem_stage_inst_dmem_ram_178__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3418) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3373 ( .A(
        mem_stage_inst_dmem_ram_178__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3419) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3372 ( .A(
        mem_stage_inst_dmem_ram_178__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3420) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3371 ( .A(
        mem_stage_inst_dmem_ram_178__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3421) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3370 ( .A(
        mem_stage_inst_dmem_ram_178__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3422) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3369 ( .A(
        mem_stage_inst_dmem_ram_178__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3423) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3368 ( .A(
        mem_stage_inst_dmem_ram_178__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3424) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3367 ( .A(
        mem_stage_inst_dmem_ram_178__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3425) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3366 ( .A(
        mem_stage_inst_dmem_ram_178__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3426) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3365 ( .A(
        mem_stage_inst_dmem_ram_178__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3427) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3364 ( .A(
        mem_stage_inst_dmem_ram_178__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5801), .Y(mem_stage_inst_dmem_n3428) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3363 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5800) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3362 ( .A(
        mem_stage_inst_dmem_ram_179__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3429) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3361 ( .A(
        mem_stage_inst_dmem_ram_179__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3430) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3360 ( .A(
        mem_stage_inst_dmem_ram_179__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3431) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3359 ( .A(
        mem_stage_inst_dmem_ram_179__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3432) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3358 ( .A(
        mem_stage_inst_dmem_ram_179__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3433) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3357 ( .A(
        mem_stage_inst_dmem_ram_179__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3434) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3356 ( .A(
        mem_stage_inst_dmem_ram_179__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3435) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3355 ( .A(
        mem_stage_inst_dmem_ram_179__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3436) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3354 ( .A(
        mem_stage_inst_dmem_ram_179__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3437) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3353 ( .A(
        mem_stage_inst_dmem_ram_179__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3438) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3352 ( .A(
        mem_stage_inst_dmem_ram_179__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3439) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3351 ( .A(
        mem_stage_inst_dmem_ram_179__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3440) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3350 ( .A(
        mem_stage_inst_dmem_ram_179__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3441) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3349 ( .A(
        mem_stage_inst_dmem_ram_179__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3442) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3348 ( .A(
        mem_stage_inst_dmem_ram_179__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3443) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3347 ( .A(
        mem_stage_inst_dmem_ram_179__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5800), .Y(mem_stage_inst_dmem_n3444) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3346 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5799) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3345 ( .A(
        mem_stage_inst_dmem_ram_180__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3445) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3344 ( .A(
        mem_stage_inst_dmem_ram_180__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3446) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3343 ( .A(
        mem_stage_inst_dmem_ram_180__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3447) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3342 ( .A(
        mem_stage_inst_dmem_ram_180__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3448) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3341 ( .A(
        mem_stage_inst_dmem_ram_180__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3449) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3340 ( .A(
        mem_stage_inst_dmem_ram_180__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3450) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3339 ( .A(
        mem_stage_inst_dmem_ram_180__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3451) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3338 ( .A(
        mem_stage_inst_dmem_ram_180__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3452) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3337 ( .A(
        mem_stage_inst_dmem_ram_180__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3453) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3336 ( .A(
        mem_stage_inst_dmem_ram_180__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3454) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3335 ( .A(
        mem_stage_inst_dmem_ram_180__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3455) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3334 ( .A(
        mem_stage_inst_dmem_ram_180__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3456) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3333 ( .A(
        mem_stage_inst_dmem_ram_180__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3457) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3332 ( .A(
        mem_stage_inst_dmem_ram_180__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3458) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3331 ( .A(
        mem_stage_inst_dmem_ram_180__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3459) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3330 ( .A(
        mem_stage_inst_dmem_ram_180__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5799), .Y(mem_stage_inst_dmem_n3460) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3329 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5798) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3328 ( .A(
        mem_stage_inst_dmem_ram_181__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3461) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3327 ( .A(
        mem_stage_inst_dmem_ram_181__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3462) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3326 ( .A(
        mem_stage_inst_dmem_ram_181__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3463) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3325 ( .A(
        mem_stage_inst_dmem_ram_181__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3464) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3324 ( .A(
        mem_stage_inst_dmem_ram_181__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3465) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3323 ( .A(
        mem_stage_inst_dmem_ram_181__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3466) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3322 ( .A(
        mem_stage_inst_dmem_ram_181__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3467) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3321 ( .A(
        mem_stage_inst_dmem_ram_181__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3468) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3320 ( .A(
        mem_stage_inst_dmem_ram_181__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3469) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3319 ( .A(
        mem_stage_inst_dmem_ram_181__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3470) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3318 ( .A(
        mem_stage_inst_dmem_ram_181__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3471) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3317 ( .A(
        mem_stage_inst_dmem_ram_181__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3472) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3316 ( .A(
        mem_stage_inst_dmem_ram_181__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3473) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3315 ( .A(
        mem_stage_inst_dmem_ram_181__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3474) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3314 ( .A(
        mem_stage_inst_dmem_ram_181__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3475) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3313 ( .A(
        mem_stage_inst_dmem_ram_181__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5798), .Y(mem_stage_inst_dmem_n3476) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3312 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5797) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3311 ( .A(
        mem_stage_inst_dmem_ram_182__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3477) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3310 ( .A(
        mem_stage_inst_dmem_ram_182__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3478) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3309 ( .A(
        mem_stage_inst_dmem_ram_182__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3479) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3308 ( .A(
        mem_stage_inst_dmem_ram_182__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3480) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3307 ( .A(
        mem_stage_inst_dmem_ram_182__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3481) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3306 ( .A(
        mem_stage_inst_dmem_ram_182__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3482) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3305 ( .A(
        mem_stage_inst_dmem_ram_182__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3483) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3304 ( .A(
        mem_stage_inst_dmem_ram_182__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3484) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3303 ( .A(
        mem_stage_inst_dmem_ram_182__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3485) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3302 ( .A(
        mem_stage_inst_dmem_ram_182__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3486) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3301 ( .A(
        mem_stage_inst_dmem_ram_182__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3487) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3300 ( .A(
        mem_stage_inst_dmem_ram_182__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3488) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3299 ( .A(
        mem_stage_inst_dmem_ram_182__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3489) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3298 ( .A(
        mem_stage_inst_dmem_ram_182__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3490) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3297 ( .A(
        mem_stage_inst_dmem_ram_182__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3491) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3296 ( .A(
        mem_stage_inst_dmem_ram_182__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5797), .Y(mem_stage_inst_dmem_n3492) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3295 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5796) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3294 ( .A(
        mem_stage_inst_dmem_ram_183__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3493) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3293 ( .A(
        mem_stage_inst_dmem_ram_183__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3494) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3292 ( .A(
        mem_stage_inst_dmem_ram_183__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3495) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3291 ( .A(
        mem_stage_inst_dmem_ram_183__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3496) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3290 ( .A(
        mem_stage_inst_dmem_ram_183__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3497) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3289 ( .A(
        mem_stage_inst_dmem_ram_183__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3498) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3288 ( .A(
        mem_stage_inst_dmem_ram_183__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3499) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3287 ( .A(
        mem_stage_inst_dmem_ram_183__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3500) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3286 ( .A(
        mem_stage_inst_dmem_ram_183__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3501) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3285 ( .A(
        mem_stage_inst_dmem_ram_183__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3502) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3284 ( .A(
        mem_stage_inst_dmem_ram_183__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3503) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3283 ( .A(
        mem_stage_inst_dmem_ram_183__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3504) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3282 ( .A(
        mem_stage_inst_dmem_ram_183__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3505) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3281 ( .A(
        mem_stage_inst_dmem_ram_183__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3506) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3280 ( .A(
        mem_stage_inst_dmem_ram_183__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3507) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3279 ( .A(
        mem_stage_inst_dmem_ram_183__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5796), .Y(mem_stage_inst_dmem_n3508) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3278 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5795) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3277 ( .A(
        mem_stage_inst_dmem_ram_184__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3509) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3276 ( .A(
        mem_stage_inst_dmem_ram_184__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3510) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3275 ( .A(
        mem_stage_inst_dmem_ram_184__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3511) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3274 ( .A(
        mem_stage_inst_dmem_ram_184__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3512) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3273 ( .A(
        mem_stage_inst_dmem_ram_184__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3513) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3272 ( .A(
        mem_stage_inst_dmem_ram_184__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3514) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3271 ( .A(
        mem_stage_inst_dmem_ram_184__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3515) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3270 ( .A(
        mem_stage_inst_dmem_ram_184__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3516) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3269 ( .A(
        mem_stage_inst_dmem_ram_184__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3517) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3268 ( .A(
        mem_stage_inst_dmem_ram_184__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3518) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3267 ( .A(
        mem_stage_inst_dmem_ram_184__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3519) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3266 ( .A(
        mem_stage_inst_dmem_ram_184__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3520) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3265 ( .A(
        mem_stage_inst_dmem_ram_184__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3521) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3264 ( .A(
        mem_stage_inst_dmem_ram_184__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3522) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3263 ( .A(
        mem_stage_inst_dmem_ram_184__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3523) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3262 ( .A(
        mem_stage_inst_dmem_ram_184__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5795), .Y(mem_stage_inst_dmem_n3524) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3261 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5794) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3260 ( .A(
        mem_stage_inst_dmem_ram_185__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3525) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3259 ( .A(
        mem_stage_inst_dmem_ram_185__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3526) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3258 ( .A(
        mem_stage_inst_dmem_ram_185__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3527) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3257 ( .A(
        mem_stage_inst_dmem_ram_185__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3528) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3256 ( .A(
        mem_stage_inst_dmem_ram_185__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3529) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3255 ( .A(
        mem_stage_inst_dmem_ram_185__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3530) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3254 ( .A(
        mem_stage_inst_dmem_ram_185__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3531) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3253 ( .A(
        mem_stage_inst_dmem_ram_185__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3532) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3252 ( .A(
        mem_stage_inst_dmem_ram_185__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3533) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3251 ( .A(
        mem_stage_inst_dmem_ram_185__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3534) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3250 ( .A(
        mem_stage_inst_dmem_ram_185__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3535) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3249 ( .A(
        mem_stage_inst_dmem_ram_185__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3536) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3248 ( .A(
        mem_stage_inst_dmem_ram_185__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3537) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3247 ( .A(
        mem_stage_inst_dmem_ram_185__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3538) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3246 ( .A(
        mem_stage_inst_dmem_ram_185__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3539) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3245 ( .A(
        mem_stage_inst_dmem_ram_185__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5794), .Y(mem_stage_inst_dmem_n3540) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3244 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5793) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3243 ( .A(
        mem_stage_inst_dmem_ram_186__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3541) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3242 ( .A(
        mem_stage_inst_dmem_ram_186__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3542) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3241 ( .A(
        mem_stage_inst_dmem_ram_186__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3543) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3240 ( .A(
        mem_stage_inst_dmem_ram_186__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3544) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3239 ( .A(
        mem_stage_inst_dmem_ram_186__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3545) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3238 ( .A(
        mem_stage_inst_dmem_ram_186__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3546) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3237 ( .A(
        mem_stage_inst_dmem_ram_186__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3547) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3236 ( .A(
        mem_stage_inst_dmem_ram_186__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3548) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3235 ( .A(
        mem_stage_inst_dmem_ram_186__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3549) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3234 ( .A(
        mem_stage_inst_dmem_ram_186__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3550) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3233 ( .A(
        mem_stage_inst_dmem_ram_186__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3551) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3232 ( .A(
        mem_stage_inst_dmem_ram_186__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3552) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3231 ( .A(
        mem_stage_inst_dmem_ram_186__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3553) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3230 ( .A(
        mem_stage_inst_dmem_ram_186__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3554) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3229 ( .A(
        mem_stage_inst_dmem_ram_186__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3555) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3228 ( .A(
        mem_stage_inst_dmem_ram_186__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5793), .Y(mem_stage_inst_dmem_n3556) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3227 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5792) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3226 ( .A(
        mem_stage_inst_dmem_ram_187__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3557) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3225 ( .A(
        mem_stage_inst_dmem_ram_187__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3558) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3224 ( .A(
        mem_stage_inst_dmem_ram_187__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3559) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3223 ( .A(
        mem_stage_inst_dmem_ram_187__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3560) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3222 ( .A(
        mem_stage_inst_dmem_ram_187__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3561) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3221 ( .A(
        mem_stage_inst_dmem_ram_187__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3562) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3220 ( .A(
        mem_stage_inst_dmem_ram_187__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3563) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3219 ( .A(
        mem_stage_inst_dmem_ram_187__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3564) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3218 ( .A(
        mem_stage_inst_dmem_ram_187__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3565) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3217 ( .A(
        mem_stage_inst_dmem_ram_187__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3566) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3216 ( .A(
        mem_stage_inst_dmem_ram_187__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3567) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3215 ( .A(
        mem_stage_inst_dmem_ram_187__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3568) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3214 ( .A(
        mem_stage_inst_dmem_ram_187__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3569) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3213 ( .A(
        mem_stage_inst_dmem_ram_187__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3570) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3212 ( .A(
        mem_stage_inst_dmem_ram_187__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3571) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3211 ( .A(
        mem_stage_inst_dmem_ram_187__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5792), .Y(mem_stage_inst_dmem_n3572) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3210 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5791) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3209 ( .A(
        mem_stage_inst_dmem_ram_188__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3573) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3208 ( .A(
        mem_stage_inst_dmem_ram_188__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3574) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3207 ( .A(
        mem_stage_inst_dmem_ram_188__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3575) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3206 ( .A(
        mem_stage_inst_dmem_ram_188__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3576) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3205 ( .A(
        mem_stage_inst_dmem_ram_188__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3577) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3204 ( .A(
        mem_stage_inst_dmem_ram_188__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3578) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3203 ( .A(
        mem_stage_inst_dmem_ram_188__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3579) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3202 ( .A(
        mem_stage_inst_dmem_ram_188__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3580) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3201 ( .A(
        mem_stage_inst_dmem_ram_188__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3581) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3200 ( .A(
        mem_stage_inst_dmem_ram_188__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3582) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3199 ( .A(
        mem_stage_inst_dmem_ram_188__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3583) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3198 ( .A(
        mem_stage_inst_dmem_ram_188__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3584) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3197 ( .A(
        mem_stage_inst_dmem_ram_188__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3585) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3196 ( .A(
        mem_stage_inst_dmem_ram_188__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3586) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3195 ( .A(
        mem_stage_inst_dmem_ram_188__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3587) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3194 ( .A(
        mem_stage_inst_dmem_ram_188__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5791), .Y(mem_stage_inst_dmem_n3588) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3193 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5790) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3192 ( .A(
        mem_stage_inst_dmem_ram_189__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3589) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3191 ( .A(
        mem_stage_inst_dmem_ram_189__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3590) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3190 ( .A(
        mem_stage_inst_dmem_ram_189__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3591) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3189 ( .A(
        mem_stage_inst_dmem_ram_189__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3592) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3188 ( .A(
        mem_stage_inst_dmem_ram_189__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3593) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3187 ( .A(
        mem_stage_inst_dmem_ram_189__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3594) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3186 ( .A(
        mem_stage_inst_dmem_ram_189__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3595) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3185 ( .A(
        mem_stage_inst_dmem_ram_189__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3596) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3184 ( .A(
        mem_stage_inst_dmem_ram_189__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3597) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3183 ( .A(
        mem_stage_inst_dmem_ram_189__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3598) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3182 ( .A(
        mem_stage_inst_dmem_ram_189__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3599) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3181 ( .A(
        mem_stage_inst_dmem_ram_189__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3600) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3180 ( .A(
        mem_stage_inst_dmem_ram_189__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3601) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3179 ( .A(
        mem_stage_inst_dmem_ram_189__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3602) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3178 ( .A(
        mem_stage_inst_dmem_ram_189__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3603) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3177 ( .A(
        mem_stage_inst_dmem_ram_189__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5790), .Y(mem_stage_inst_dmem_n3604) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3176 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5789) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3175 ( .A(
        mem_stage_inst_dmem_ram_190__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3605) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3174 ( .A(
        mem_stage_inst_dmem_ram_190__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3606) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3173 ( .A(
        mem_stage_inst_dmem_ram_190__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3607) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3172 ( .A(
        mem_stage_inst_dmem_ram_190__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3608) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3171 ( .A(
        mem_stage_inst_dmem_ram_190__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3609) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3170 ( .A(
        mem_stage_inst_dmem_ram_190__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3610) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3169 ( .A(
        mem_stage_inst_dmem_ram_190__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3611) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3168 ( .A(
        mem_stage_inst_dmem_ram_190__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3612) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3167 ( .A(
        mem_stage_inst_dmem_ram_190__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3613) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3166 ( .A(
        mem_stage_inst_dmem_ram_190__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3614) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3165 ( .A(
        mem_stage_inst_dmem_ram_190__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3615) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3164 ( .A(
        mem_stage_inst_dmem_ram_190__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3616) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3163 ( .A(
        mem_stage_inst_dmem_ram_190__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3617) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3162 ( .A(
        mem_stage_inst_dmem_ram_190__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3618) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3161 ( .A(
        mem_stage_inst_dmem_ram_190__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3619) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3160 ( .A(
        mem_stage_inst_dmem_ram_190__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5789), .Y(mem_stage_inst_dmem_n3620) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3159 ( .A(mem_stage_inst_dmem_n5788), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5787) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3158 ( .A(
        mem_stage_inst_dmem_ram_191__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3621) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3157 ( .A(
        mem_stage_inst_dmem_ram_191__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3622) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3156 ( .A(
        mem_stage_inst_dmem_ram_191__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3623) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3155 ( .A(
        mem_stage_inst_dmem_ram_191__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3624) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3154 ( .A(
        mem_stage_inst_dmem_ram_191__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3625) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3153 ( .A(
        mem_stage_inst_dmem_ram_191__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3626) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3152 ( .A(
        mem_stage_inst_dmem_ram_191__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3627) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3151 ( .A(
        mem_stage_inst_dmem_ram_191__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3628) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3150 ( .A(
        mem_stage_inst_dmem_ram_191__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3629) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3149 ( .A(
        mem_stage_inst_dmem_ram_191__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3630) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3148 ( .A(
        mem_stage_inst_dmem_ram_191__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3631) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3147 ( .A(
        mem_stage_inst_dmem_ram_191__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3632) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3146 ( .A(
        mem_stage_inst_dmem_ram_191__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3633) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3145 ( .A(
        mem_stage_inst_dmem_ram_191__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3634) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3144 ( .A(
        mem_stage_inst_dmem_ram_191__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3635) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3143 ( .A(
        mem_stage_inst_dmem_ram_191__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5787), .Y(mem_stage_inst_dmem_n3636) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3142 ( .A(mem_stage_inst_dmem_n5786), 
        .B(ex_pipeline_reg_out[28]), .Y(mem_stage_inst_dmem_n5731) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3141 ( .A(mem_stage_inst_dmem_n5731), 
        .B(mem_stage_inst_dmem_n5712), .Y(mem_stage_inst_dmem_n5770) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3140 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5785) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3139 ( .A(
        mem_stage_inst_dmem_ram_192__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3637) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3138 ( .A(
        mem_stage_inst_dmem_ram_192__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3638) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3137 ( .A(
        mem_stage_inst_dmem_ram_192__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3639) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3136 ( .A(
        mem_stage_inst_dmem_ram_192__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3640) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3135 ( .A(
        mem_stage_inst_dmem_ram_192__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3641) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3134 ( .A(
        mem_stage_inst_dmem_ram_192__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3642) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3133 ( .A(
        mem_stage_inst_dmem_ram_192__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3643) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3132 ( .A(
        mem_stage_inst_dmem_ram_192__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3644) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3131 ( .A(
        mem_stage_inst_dmem_ram_192__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3645) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3130 ( .A(
        mem_stage_inst_dmem_ram_192__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3646) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3129 ( .A(
        mem_stage_inst_dmem_ram_192__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3647) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3128 ( .A(
        mem_stage_inst_dmem_ram_192__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3648) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3127 ( .A(
        mem_stage_inst_dmem_ram_192__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3649) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3126 ( .A(
        mem_stage_inst_dmem_ram_192__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3650) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3125 ( .A(
        mem_stage_inst_dmem_ram_192__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3651) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3124 ( .A(
        mem_stage_inst_dmem_ram_192__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5785), .Y(mem_stage_inst_dmem_n3652) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3123 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5784) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3122 ( .A(
        mem_stage_inst_dmem_ram_193__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3653) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3121 ( .A(
        mem_stage_inst_dmem_ram_193__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3654) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3120 ( .A(
        mem_stage_inst_dmem_ram_193__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3655) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3119 ( .A(
        mem_stage_inst_dmem_ram_193__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3656) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3118 ( .A(
        mem_stage_inst_dmem_ram_193__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3657) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3117 ( .A(
        mem_stage_inst_dmem_ram_193__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3658) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3116 ( .A(
        mem_stage_inst_dmem_ram_193__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3659) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3115 ( .A(
        mem_stage_inst_dmem_ram_193__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3660) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3114 ( .A(
        mem_stage_inst_dmem_ram_193__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3661) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3113 ( .A(
        mem_stage_inst_dmem_ram_193__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3662) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3112 ( .A(
        mem_stage_inst_dmem_ram_193__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3663) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3111 ( .A(
        mem_stage_inst_dmem_ram_193__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3664) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3110 ( .A(
        mem_stage_inst_dmem_ram_193__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3665) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3109 ( .A(
        mem_stage_inst_dmem_ram_193__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3666) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3108 ( .A(
        mem_stage_inst_dmem_ram_193__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3667) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3107 ( .A(
        mem_stage_inst_dmem_ram_193__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5784), .Y(mem_stage_inst_dmem_n3668) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3106 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5783) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3105 ( .A(
        mem_stage_inst_dmem_ram_194__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3669) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3104 ( .A(
        mem_stage_inst_dmem_ram_194__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3670) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3103 ( .A(
        mem_stage_inst_dmem_ram_194__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3671) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3102 ( .A(
        mem_stage_inst_dmem_ram_194__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3672) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3101 ( .A(
        mem_stage_inst_dmem_ram_194__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3673) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3100 ( .A(
        mem_stage_inst_dmem_ram_194__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3674) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3099 ( .A(
        mem_stage_inst_dmem_ram_194__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3675) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3098 ( .A(
        mem_stage_inst_dmem_ram_194__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3676) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3097 ( .A(
        mem_stage_inst_dmem_ram_194__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3677) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3096 ( .A(
        mem_stage_inst_dmem_ram_194__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3678) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3095 ( .A(
        mem_stage_inst_dmem_ram_194__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3679) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3094 ( .A(
        mem_stage_inst_dmem_ram_194__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3680) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3093 ( .A(
        mem_stage_inst_dmem_ram_194__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3681) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3092 ( .A(
        mem_stage_inst_dmem_ram_194__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3682) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3091 ( .A(
        mem_stage_inst_dmem_ram_194__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3683) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3090 ( .A(
        mem_stage_inst_dmem_ram_194__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5783), .Y(mem_stage_inst_dmem_n3684) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3089 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5782) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3088 ( .A(
        mem_stage_inst_dmem_ram_195__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3685) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3087 ( .A(
        mem_stage_inst_dmem_ram_195__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3686) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3086 ( .A(
        mem_stage_inst_dmem_ram_195__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3687) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3085 ( .A(
        mem_stage_inst_dmem_ram_195__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3688) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3084 ( .A(
        mem_stage_inst_dmem_ram_195__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3689) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3083 ( .A(
        mem_stage_inst_dmem_ram_195__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3690) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3082 ( .A(
        mem_stage_inst_dmem_ram_195__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3691) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3081 ( .A(
        mem_stage_inst_dmem_ram_195__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3692) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3080 ( .A(
        mem_stage_inst_dmem_ram_195__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3693) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3079 ( .A(
        mem_stage_inst_dmem_ram_195__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3694) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3078 ( .A(
        mem_stage_inst_dmem_ram_195__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3695) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3077 ( .A(
        mem_stage_inst_dmem_ram_195__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3696) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3076 ( .A(
        mem_stage_inst_dmem_ram_195__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3697) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3075 ( .A(
        mem_stage_inst_dmem_ram_195__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3698) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3074 ( .A(
        mem_stage_inst_dmem_ram_195__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3699) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3073 ( .A(
        mem_stage_inst_dmem_ram_195__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5782), .Y(mem_stage_inst_dmem_n3700) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3072 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5781) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3071 ( .A(
        mem_stage_inst_dmem_ram_196__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3701) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3070 ( .A(
        mem_stage_inst_dmem_ram_196__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3702) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3069 ( .A(
        mem_stage_inst_dmem_ram_196__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3703) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3068 ( .A(
        mem_stage_inst_dmem_ram_196__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3704) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3067 ( .A(
        mem_stage_inst_dmem_ram_196__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3705) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3066 ( .A(
        mem_stage_inst_dmem_ram_196__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3706) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3065 ( .A(
        mem_stage_inst_dmem_ram_196__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3707) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3064 ( .A(
        mem_stage_inst_dmem_ram_196__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3708) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3063 ( .A(
        mem_stage_inst_dmem_ram_196__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3709) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3062 ( .A(
        mem_stage_inst_dmem_ram_196__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3710) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3061 ( .A(
        mem_stage_inst_dmem_ram_196__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3711) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3060 ( .A(
        mem_stage_inst_dmem_ram_196__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3712) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3059 ( .A(
        mem_stage_inst_dmem_ram_196__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3713) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3058 ( .A(
        mem_stage_inst_dmem_ram_196__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3714) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3057 ( .A(
        mem_stage_inst_dmem_ram_196__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3715) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3056 ( .A(
        mem_stage_inst_dmem_ram_196__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5781), .Y(mem_stage_inst_dmem_n3716) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3055 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5780) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3054 ( .A(
        mem_stage_inst_dmem_ram_197__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3717) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3053 ( .A(
        mem_stage_inst_dmem_ram_197__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3718) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3052 ( .A(
        mem_stage_inst_dmem_ram_197__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3719) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3051 ( .A(
        mem_stage_inst_dmem_ram_197__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3720) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3050 ( .A(
        mem_stage_inst_dmem_ram_197__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3721) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3049 ( .A(
        mem_stage_inst_dmem_ram_197__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3722) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3048 ( .A(
        mem_stage_inst_dmem_ram_197__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3723) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3047 ( .A(
        mem_stage_inst_dmem_ram_197__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3724) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3046 ( .A(
        mem_stage_inst_dmem_ram_197__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3725) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3045 ( .A(
        mem_stage_inst_dmem_ram_197__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3726) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3044 ( .A(
        mem_stage_inst_dmem_ram_197__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3727) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3043 ( .A(
        mem_stage_inst_dmem_ram_197__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3728) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3042 ( .A(
        mem_stage_inst_dmem_ram_197__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3729) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3041 ( .A(
        mem_stage_inst_dmem_ram_197__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3730) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3040 ( .A(
        mem_stage_inst_dmem_ram_197__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3731) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3039 ( .A(
        mem_stage_inst_dmem_ram_197__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5780), .Y(mem_stage_inst_dmem_n3732) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3038 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5779) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3037 ( .A(
        mem_stage_inst_dmem_ram_198__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3733) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3036 ( .A(
        mem_stage_inst_dmem_ram_198__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3734) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3035 ( .A(
        mem_stage_inst_dmem_ram_198__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3735) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3034 ( .A(
        mem_stage_inst_dmem_ram_198__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3736) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3033 ( .A(
        mem_stage_inst_dmem_ram_198__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3737) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3032 ( .A(
        mem_stage_inst_dmem_ram_198__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3738) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3031 ( .A(
        mem_stage_inst_dmem_ram_198__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3739) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3030 ( .A(
        mem_stage_inst_dmem_ram_198__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3740) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3029 ( .A(
        mem_stage_inst_dmem_ram_198__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3741) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3028 ( .A(
        mem_stage_inst_dmem_ram_198__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3742) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3027 ( .A(
        mem_stage_inst_dmem_ram_198__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3743) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3026 ( .A(
        mem_stage_inst_dmem_ram_198__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3744) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3025 ( .A(
        mem_stage_inst_dmem_ram_198__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3745) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3024 ( .A(
        mem_stage_inst_dmem_ram_198__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3746) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3023 ( .A(
        mem_stage_inst_dmem_ram_198__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3747) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3022 ( .A(
        mem_stage_inst_dmem_ram_198__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5779), .Y(mem_stage_inst_dmem_n3748) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3021 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5778) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3020 ( .A(
        mem_stage_inst_dmem_ram_199__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3749) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3019 ( .A(
        mem_stage_inst_dmem_ram_199__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3750) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3018 ( .A(
        mem_stage_inst_dmem_ram_199__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3751) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3017 ( .A(
        mem_stage_inst_dmem_ram_199__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3752) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3016 ( .A(
        mem_stage_inst_dmem_ram_199__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3753) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3015 ( .A(
        mem_stage_inst_dmem_ram_199__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3754) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3014 ( .A(
        mem_stage_inst_dmem_ram_199__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3755) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3013 ( .A(
        mem_stage_inst_dmem_ram_199__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3756) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3012 ( .A(
        mem_stage_inst_dmem_ram_199__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3757) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3011 ( .A(
        mem_stage_inst_dmem_ram_199__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3758) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3010 ( .A(
        mem_stage_inst_dmem_ram_199__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3759) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3009 ( .A(
        mem_stage_inst_dmem_ram_199__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3760) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3008 ( .A(
        mem_stage_inst_dmem_ram_199__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3761) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3007 ( .A(
        mem_stage_inst_dmem_ram_199__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3762) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3006 ( .A(
        mem_stage_inst_dmem_ram_199__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3763) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3005 ( .A(
        mem_stage_inst_dmem_ram_199__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5778), .Y(mem_stage_inst_dmem_n3764) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u3004 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5777) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3003 ( .A(
        mem_stage_inst_dmem_ram_200__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3765) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3002 ( .A(
        mem_stage_inst_dmem_ram_200__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3766) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3001 ( .A(
        mem_stage_inst_dmem_ram_200__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3767) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u3000 ( .A(
        mem_stage_inst_dmem_ram_200__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3768) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2999 ( .A(
        mem_stage_inst_dmem_ram_200__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3769) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2998 ( .A(
        mem_stage_inst_dmem_ram_200__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3770) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2997 ( .A(
        mem_stage_inst_dmem_ram_200__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3771) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2996 ( .A(
        mem_stage_inst_dmem_ram_200__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3772) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2995 ( .A(
        mem_stage_inst_dmem_ram_200__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3773) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2994 ( .A(
        mem_stage_inst_dmem_ram_200__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3774) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2993 ( .A(
        mem_stage_inst_dmem_ram_200__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3775) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2992 ( .A(
        mem_stage_inst_dmem_ram_200__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3776) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2991 ( .A(
        mem_stage_inst_dmem_ram_200__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3777) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2990 ( .A(
        mem_stage_inst_dmem_ram_200__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3778) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2989 ( .A(
        mem_stage_inst_dmem_ram_200__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3779) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2988 ( .A(
        mem_stage_inst_dmem_ram_200__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5777), .Y(mem_stage_inst_dmem_n3780) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2987 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5776) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2986 ( .A(
        mem_stage_inst_dmem_ram_201__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3781) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2985 ( .A(
        mem_stage_inst_dmem_ram_201__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3782) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2984 ( .A(
        mem_stage_inst_dmem_ram_201__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3783) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2983 ( .A(
        mem_stage_inst_dmem_ram_201__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3784) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2982 ( .A(
        mem_stage_inst_dmem_ram_201__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3785) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2981 ( .A(
        mem_stage_inst_dmem_ram_201__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3786) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2980 ( .A(
        mem_stage_inst_dmem_ram_201__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3787) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2979 ( .A(
        mem_stage_inst_dmem_ram_201__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3788) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2978 ( .A(
        mem_stage_inst_dmem_ram_201__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3789) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2977 ( .A(
        mem_stage_inst_dmem_ram_201__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3790) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2976 ( .A(
        mem_stage_inst_dmem_ram_201__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3791) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2975 ( .A(
        mem_stage_inst_dmem_ram_201__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3792) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2974 ( .A(
        mem_stage_inst_dmem_ram_201__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3793) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2973 ( .A(
        mem_stage_inst_dmem_ram_201__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3794) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2972 ( .A(
        mem_stage_inst_dmem_ram_201__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3795) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2971 ( .A(
        mem_stage_inst_dmem_ram_201__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5776), .Y(mem_stage_inst_dmem_n3796) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2970 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5775) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2969 ( .A(
        mem_stage_inst_dmem_ram_202__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3797) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2968 ( .A(
        mem_stage_inst_dmem_ram_202__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3798) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2967 ( .A(
        mem_stage_inst_dmem_ram_202__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3799) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2966 ( .A(
        mem_stage_inst_dmem_ram_202__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3800) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2965 ( .A(
        mem_stage_inst_dmem_ram_202__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3801) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2964 ( .A(
        mem_stage_inst_dmem_ram_202__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3802) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2963 ( .A(
        mem_stage_inst_dmem_ram_202__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3803) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2962 ( .A(
        mem_stage_inst_dmem_ram_202__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3804) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2961 ( .A(
        mem_stage_inst_dmem_ram_202__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3805) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2960 ( .A(
        mem_stage_inst_dmem_ram_202__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3806) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2959 ( .A(
        mem_stage_inst_dmem_ram_202__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3807) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2958 ( .A(
        mem_stage_inst_dmem_ram_202__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3808) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2957 ( .A(
        mem_stage_inst_dmem_ram_202__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3809) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2956 ( .A(
        mem_stage_inst_dmem_ram_202__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3810) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2955 ( .A(
        mem_stage_inst_dmem_ram_202__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3811) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2954 ( .A(
        mem_stage_inst_dmem_ram_202__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5775), .Y(mem_stage_inst_dmem_n3812) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2953 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5774) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2952 ( .A(
        mem_stage_inst_dmem_ram_203__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3813) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2951 ( .A(
        mem_stage_inst_dmem_ram_203__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3814) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2950 ( .A(
        mem_stage_inst_dmem_ram_203__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3815) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2949 ( .A(
        mem_stage_inst_dmem_ram_203__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3816) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2948 ( .A(
        mem_stage_inst_dmem_ram_203__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3817) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2947 ( .A(
        mem_stage_inst_dmem_ram_203__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3818) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2946 ( .A(
        mem_stage_inst_dmem_ram_203__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3819) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2945 ( .A(
        mem_stage_inst_dmem_ram_203__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3820) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2944 ( .A(
        mem_stage_inst_dmem_ram_203__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3821) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2943 ( .A(
        mem_stage_inst_dmem_ram_203__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3822) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2942 ( .A(
        mem_stage_inst_dmem_ram_203__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3823) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2941 ( .A(
        mem_stage_inst_dmem_ram_203__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3824) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2940 ( .A(
        mem_stage_inst_dmem_ram_203__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3825) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2939 ( .A(
        mem_stage_inst_dmem_ram_203__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3826) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2938 ( .A(
        mem_stage_inst_dmem_ram_203__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3827) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2937 ( .A(
        mem_stage_inst_dmem_ram_203__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5774), .Y(mem_stage_inst_dmem_n3828) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2936 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5773) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2935 ( .A(
        mem_stage_inst_dmem_ram_204__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3829) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2934 ( .A(
        mem_stage_inst_dmem_ram_204__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3830) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2933 ( .A(
        mem_stage_inst_dmem_ram_204__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3831) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2932 ( .A(
        mem_stage_inst_dmem_ram_204__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3832) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2931 ( .A(
        mem_stage_inst_dmem_ram_204__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3833) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2930 ( .A(
        mem_stage_inst_dmem_ram_204__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3834) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2929 ( .A(
        mem_stage_inst_dmem_ram_204__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3835) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2928 ( .A(
        mem_stage_inst_dmem_ram_204__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3836) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2927 ( .A(
        mem_stage_inst_dmem_ram_204__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3837) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2926 ( .A(
        mem_stage_inst_dmem_ram_204__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3838) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2925 ( .A(
        mem_stage_inst_dmem_ram_204__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3839) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2924 ( .A(
        mem_stage_inst_dmem_ram_204__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3840) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2923 ( .A(
        mem_stage_inst_dmem_ram_204__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3841) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2922 ( .A(
        mem_stage_inst_dmem_ram_204__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3842) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2921 ( .A(
        mem_stage_inst_dmem_ram_204__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3843) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2920 ( .A(
        mem_stage_inst_dmem_ram_204__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5773), .Y(mem_stage_inst_dmem_n3844) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2919 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5772) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2918 ( .A(
        mem_stage_inst_dmem_ram_205__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3845) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2917 ( .A(
        mem_stage_inst_dmem_ram_205__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3846) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2916 ( .A(
        mem_stage_inst_dmem_ram_205__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3847) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2915 ( .A(
        mem_stage_inst_dmem_ram_205__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3848) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2914 ( .A(
        mem_stage_inst_dmem_ram_205__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3849) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2913 ( .A(
        mem_stage_inst_dmem_ram_205__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3850) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2912 ( .A(
        mem_stage_inst_dmem_ram_205__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3851) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2911 ( .A(
        mem_stage_inst_dmem_ram_205__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3852) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2910 ( .A(
        mem_stage_inst_dmem_ram_205__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3853) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2909 ( .A(
        mem_stage_inst_dmem_ram_205__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3854) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2908 ( .A(
        mem_stage_inst_dmem_ram_205__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3855) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2907 ( .A(
        mem_stage_inst_dmem_ram_205__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3856) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2906 ( .A(
        mem_stage_inst_dmem_ram_205__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3857) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2905 ( .A(
        mem_stage_inst_dmem_ram_205__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3858) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2904 ( .A(
        mem_stage_inst_dmem_ram_205__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3859) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2903 ( .A(
        mem_stage_inst_dmem_ram_205__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5772), .Y(mem_stage_inst_dmem_n3860) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2902 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5771) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2901 ( .A(
        mem_stage_inst_dmem_ram_206__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3861) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2900 ( .A(
        mem_stage_inst_dmem_ram_206__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3862) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2899 ( .A(
        mem_stage_inst_dmem_ram_206__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3863) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2898 ( .A(
        mem_stage_inst_dmem_ram_206__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3864) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2897 ( .A(
        mem_stage_inst_dmem_ram_206__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3865) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2896 ( .A(
        mem_stage_inst_dmem_ram_206__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3866) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2895 ( .A(
        mem_stage_inst_dmem_ram_206__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3867) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2894 ( .A(
        mem_stage_inst_dmem_ram_206__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3868) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2893 ( .A(
        mem_stage_inst_dmem_ram_206__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3869) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2892 ( .A(
        mem_stage_inst_dmem_ram_206__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3870) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2891 ( .A(
        mem_stage_inst_dmem_ram_206__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3871) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2890 ( .A(
        mem_stage_inst_dmem_ram_206__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3872) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2889 ( .A(
        mem_stage_inst_dmem_ram_206__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3873) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2888 ( .A(
        mem_stage_inst_dmem_ram_206__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3874) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2887 ( .A(
        mem_stage_inst_dmem_ram_206__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3875) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2886 ( .A(
        mem_stage_inst_dmem_ram_206__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5771), .Y(mem_stage_inst_dmem_n3876) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2885 ( .A(mem_stage_inst_dmem_n5770), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5769) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2884 ( .A(
        mem_stage_inst_dmem_ram_207__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3877) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2883 ( .A(
        mem_stage_inst_dmem_ram_207__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3878) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2882 ( .A(
        mem_stage_inst_dmem_ram_207__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3879) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2881 ( .A(
        mem_stage_inst_dmem_ram_207__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3880) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2880 ( .A(
        mem_stage_inst_dmem_ram_207__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3881) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2879 ( .A(
        mem_stage_inst_dmem_ram_207__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3882) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2878 ( .A(
        mem_stage_inst_dmem_ram_207__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3883) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2877 ( .A(
        mem_stage_inst_dmem_ram_207__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3884) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2876 ( .A(
        mem_stage_inst_dmem_ram_207__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3885) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2875 ( .A(
        mem_stage_inst_dmem_ram_207__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3886) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2874 ( .A(
        mem_stage_inst_dmem_ram_207__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3887) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2873 ( .A(
        mem_stage_inst_dmem_ram_207__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3888) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2872 ( .A(
        mem_stage_inst_dmem_ram_207__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3889) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2871 ( .A(
        mem_stage_inst_dmem_ram_207__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3890) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2870 ( .A(
        mem_stage_inst_dmem_ram_207__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3891) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2869 ( .A(
        mem_stage_inst_dmem_ram_207__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5769), .Y(mem_stage_inst_dmem_n3892) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2868 ( .A(mem_stage_inst_dmem_n5731), 
        .B(mem_stage_inst_dmem_n5768), .Y(mem_stage_inst_dmem_n5752) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2867 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5767) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2866 ( .A(
        mem_stage_inst_dmem_ram_208__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3893) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2865 ( .A(
        mem_stage_inst_dmem_ram_208__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3894) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2864 ( .A(
        mem_stage_inst_dmem_ram_208__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3895) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2863 ( .A(
        mem_stage_inst_dmem_ram_208__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3896) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2862 ( .A(
        mem_stage_inst_dmem_ram_208__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3897) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2861 ( .A(
        mem_stage_inst_dmem_ram_208__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3898) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2860 ( .A(
        mem_stage_inst_dmem_ram_208__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3899) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2859 ( .A(
        mem_stage_inst_dmem_ram_208__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3900) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2858 ( .A(
        mem_stage_inst_dmem_ram_208__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3901) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2857 ( .A(
        mem_stage_inst_dmem_ram_208__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3902) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2856 ( .A(
        mem_stage_inst_dmem_ram_208__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3903) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2855 ( .A(
        mem_stage_inst_dmem_ram_208__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3904) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2854 ( .A(
        mem_stage_inst_dmem_ram_208__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3905) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2853 ( .A(
        mem_stage_inst_dmem_ram_208__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3906) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2852 ( .A(
        mem_stage_inst_dmem_ram_208__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3907) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2851 ( .A(
        mem_stage_inst_dmem_ram_208__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5767), .Y(mem_stage_inst_dmem_n3908) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2850 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5766) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2849 ( .A(
        mem_stage_inst_dmem_ram_209__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3909) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2848 ( .A(
        mem_stage_inst_dmem_ram_209__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3910) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2847 ( .A(
        mem_stage_inst_dmem_ram_209__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3911) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2846 ( .A(
        mem_stage_inst_dmem_ram_209__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3912) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2845 ( .A(
        mem_stage_inst_dmem_ram_209__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3913) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2844 ( .A(
        mem_stage_inst_dmem_ram_209__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3914) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2843 ( .A(
        mem_stage_inst_dmem_ram_209__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3915) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2842 ( .A(
        mem_stage_inst_dmem_ram_209__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3916) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2841 ( .A(
        mem_stage_inst_dmem_ram_209__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3917) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2840 ( .A(
        mem_stage_inst_dmem_ram_209__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3918) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2839 ( .A(
        mem_stage_inst_dmem_ram_209__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3919) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2838 ( .A(
        mem_stage_inst_dmem_ram_209__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3920) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2837 ( .A(
        mem_stage_inst_dmem_ram_209__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3921) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2836 ( .A(
        mem_stage_inst_dmem_ram_209__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3922) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2835 ( .A(
        mem_stage_inst_dmem_ram_209__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3923) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2834 ( .A(
        mem_stage_inst_dmem_ram_209__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5766), .Y(mem_stage_inst_dmem_n3924) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2833 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5765) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2832 ( .A(
        mem_stage_inst_dmem_ram_210__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3925) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2831 ( .A(
        mem_stage_inst_dmem_ram_210__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3926) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2830 ( .A(
        mem_stage_inst_dmem_ram_210__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3927) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2829 ( .A(
        mem_stage_inst_dmem_ram_210__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3928) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2828 ( .A(
        mem_stage_inst_dmem_ram_210__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3929) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2827 ( .A(
        mem_stage_inst_dmem_ram_210__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3930) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2826 ( .A(
        mem_stage_inst_dmem_ram_210__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3931) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2825 ( .A(
        mem_stage_inst_dmem_ram_210__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3932) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2824 ( .A(
        mem_stage_inst_dmem_ram_210__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3933) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2823 ( .A(
        mem_stage_inst_dmem_ram_210__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3934) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2822 ( .A(
        mem_stage_inst_dmem_ram_210__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3935) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2821 ( .A(
        mem_stage_inst_dmem_ram_210__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3936) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2820 ( .A(
        mem_stage_inst_dmem_ram_210__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3937) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2819 ( .A(
        mem_stage_inst_dmem_ram_210__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3938) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2818 ( .A(
        mem_stage_inst_dmem_ram_210__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3939) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2817 ( .A(
        mem_stage_inst_dmem_ram_210__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5765), .Y(mem_stage_inst_dmem_n3940) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2816 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5764) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2815 ( .A(
        mem_stage_inst_dmem_ram_211__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3941) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2814 ( .A(
        mem_stage_inst_dmem_ram_211__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3942) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2813 ( .A(
        mem_stage_inst_dmem_ram_211__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3943) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2812 ( .A(
        mem_stage_inst_dmem_ram_211__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3944) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2811 ( .A(
        mem_stage_inst_dmem_ram_211__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3945) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2810 ( .A(
        mem_stage_inst_dmem_ram_211__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3946) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2809 ( .A(
        mem_stage_inst_dmem_ram_211__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3947) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2808 ( .A(
        mem_stage_inst_dmem_ram_211__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3948) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2807 ( .A(
        mem_stage_inst_dmem_ram_211__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3949) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2806 ( .A(
        mem_stage_inst_dmem_ram_211__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3950) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2805 ( .A(
        mem_stage_inst_dmem_ram_211__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3951) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2804 ( .A(
        mem_stage_inst_dmem_ram_211__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3952) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2803 ( .A(
        mem_stage_inst_dmem_ram_211__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3953) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2802 ( .A(
        mem_stage_inst_dmem_ram_211__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3954) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2801 ( .A(
        mem_stage_inst_dmem_ram_211__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3955) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2800 ( .A(
        mem_stage_inst_dmem_ram_211__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5764), .Y(mem_stage_inst_dmem_n3956) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2799 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5763) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2798 ( .A(
        mem_stage_inst_dmem_ram_212__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3957) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2797 ( .A(
        mem_stage_inst_dmem_ram_212__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3958) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2796 ( .A(
        mem_stage_inst_dmem_ram_212__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3959) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2795 ( .A(
        mem_stage_inst_dmem_ram_212__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3960) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2794 ( .A(
        mem_stage_inst_dmem_ram_212__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3961) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2793 ( .A(
        mem_stage_inst_dmem_ram_212__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3962) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2792 ( .A(
        mem_stage_inst_dmem_ram_212__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3963) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2791 ( .A(
        mem_stage_inst_dmem_ram_212__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3964) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2790 ( .A(
        mem_stage_inst_dmem_ram_212__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3965) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2789 ( .A(
        mem_stage_inst_dmem_ram_212__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3966) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2788 ( .A(
        mem_stage_inst_dmem_ram_212__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3967) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2787 ( .A(
        mem_stage_inst_dmem_ram_212__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3968) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2786 ( .A(
        mem_stage_inst_dmem_ram_212__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3969) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2785 ( .A(
        mem_stage_inst_dmem_ram_212__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3970) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2784 ( .A(
        mem_stage_inst_dmem_ram_212__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3971) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2783 ( .A(
        mem_stage_inst_dmem_ram_212__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5763), .Y(mem_stage_inst_dmem_n3972) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2782 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5762) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2781 ( .A(
        mem_stage_inst_dmem_ram_213__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3973) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2780 ( .A(
        mem_stage_inst_dmem_ram_213__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3974) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2779 ( .A(
        mem_stage_inst_dmem_ram_213__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3975) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2778 ( .A(
        mem_stage_inst_dmem_ram_213__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3976) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2777 ( .A(
        mem_stage_inst_dmem_ram_213__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3977) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2776 ( .A(
        mem_stage_inst_dmem_ram_213__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3978) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2775 ( .A(
        mem_stage_inst_dmem_ram_213__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3979) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2774 ( .A(
        mem_stage_inst_dmem_ram_213__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3980) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2773 ( .A(
        mem_stage_inst_dmem_ram_213__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3981) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2772 ( .A(
        mem_stage_inst_dmem_ram_213__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3982) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2771 ( .A(
        mem_stage_inst_dmem_ram_213__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3983) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2770 ( .A(
        mem_stage_inst_dmem_ram_213__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3984) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2769 ( .A(
        mem_stage_inst_dmem_ram_213__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3985) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2768 ( .A(
        mem_stage_inst_dmem_ram_213__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3986) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2767 ( .A(
        mem_stage_inst_dmem_ram_213__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3987) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2766 ( .A(
        mem_stage_inst_dmem_ram_213__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5762), .Y(mem_stage_inst_dmem_n3988) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2765 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5761) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2764 ( .A(
        mem_stage_inst_dmem_ram_214__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3989) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2763 ( .A(
        mem_stage_inst_dmem_ram_214__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3990) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2762 ( .A(
        mem_stage_inst_dmem_ram_214__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3991) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2761 ( .A(
        mem_stage_inst_dmem_ram_214__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3992) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2760 ( .A(
        mem_stage_inst_dmem_ram_214__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3993) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2759 ( .A(
        mem_stage_inst_dmem_ram_214__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3994) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2758 ( .A(
        mem_stage_inst_dmem_ram_214__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3995) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2757 ( .A(
        mem_stage_inst_dmem_ram_214__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3996) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2756 ( .A(
        mem_stage_inst_dmem_ram_214__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3997) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2755 ( .A(
        mem_stage_inst_dmem_ram_214__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3998) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2754 ( .A(
        mem_stage_inst_dmem_ram_214__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n3999) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2753 ( .A(
        mem_stage_inst_dmem_ram_214__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n4000) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2752 ( .A(
        mem_stage_inst_dmem_ram_214__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n4001) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2751 ( .A(
        mem_stage_inst_dmem_ram_214__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n4002) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2750 ( .A(
        mem_stage_inst_dmem_ram_214__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n4003) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2749 ( .A(
        mem_stage_inst_dmem_ram_214__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5761), .Y(mem_stage_inst_dmem_n4004) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2748 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5760) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2747 ( .A(
        mem_stage_inst_dmem_ram_215__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4005) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2746 ( .A(
        mem_stage_inst_dmem_ram_215__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4006) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2745 ( .A(
        mem_stage_inst_dmem_ram_215__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4007) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2744 ( .A(
        mem_stage_inst_dmem_ram_215__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4008) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2743 ( .A(
        mem_stage_inst_dmem_ram_215__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4009) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2742 ( .A(
        mem_stage_inst_dmem_ram_215__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4010) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2741 ( .A(
        mem_stage_inst_dmem_ram_215__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4011) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2740 ( .A(
        mem_stage_inst_dmem_ram_215__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4012) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2739 ( .A(
        mem_stage_inst_dmem_ram_215__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4013) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2738 ( .A(
        mem_stage_inst_dmem_ram_215__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4014) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2737 ( .A(
        mem_stage_inst_dmem_ram_215__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4015) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2736 ( .A(
        mem_stage_inst_dmem_ram_215__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4016) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2735 ( .A(
        mem_stage_inst_dmem_ram_215__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4017) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2734 ( .A(
        mem_stage_inst_dmem_ram_215__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4018) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2733 ( .A(
        mem_stage_inst_dmem_ram_215__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4019) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2732 ( .A(
        mem_stage_inst_dmem_ram_215__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5760), .Y(mem_stage_inst_dmem_n4020) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2731 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5759) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2730 ( .A(
        mem_stage_inst_dmem_ram_216__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4021) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2729 ( .A(
        mem_stage_inst_dmem_ram_216__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4022) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2728 ( .A(
        mem_stage_inst_dmem_ram_216__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4023) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2727 ( .A(
        mem_stage_inst_dmem_ram_216__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4024) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2726 ( .A(
        mem_stage_inst_dmem_ram_216__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4025) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2725 ( .A(
        mem_stage_inst_dmem_ram_216__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4026) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2724 ( .A(
        mem_stage_inst_dmem_ram_216__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4027) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2723 ( .A(
        mem_stage_inst_dmem_ram_216__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4028) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2722 ( .A(
        mem_stage_inst_dmem_ram_216__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4029) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2721 ( .A(
        mem_stage_inst_dmem_ram_216__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4030) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2720 ( .A(
        mem_stage_inst_dmem_ram_216__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4031) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2719 ( .A(
        mem_stage_inst_dmem_ram_216__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4032) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2718 ( .A(
        mem_stage_inst_dmem_ram_216__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4033) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2717 ( .A(
        mem_stage_inst_dmem_ram_216__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4034) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2716 ( .A(
        mem_stage_inst_dmem_ram_216__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4035) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2715 ( .A(
        mem_stage_inst_dmem_ram_216__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5759), .Y(mem_stage_inst_dmem_n4036) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2714 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5758) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2713 ( .A(
        mem_stage_inst_dmem_ram_217__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4037) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2712 ( .A(
        mem_stage_inst_dmem_ram_217__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4038) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2711 ( .A(
        mem_stage_inst_dmem_ram_217__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4039) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2710 ( .A(
        mem_stage_inst_dmem_ram_217__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4040) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2709 ( .A(
        mem_stage_inst_dmem_ram_217__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4041) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2708 ( .A(
        mem_stage_inst_dmem_ram_217__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4042) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2707 ( .A(
        mem_stage_inst_dmem_ram_217__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4043) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2706 ( .A(
        mem_stage_inst_dmem_ram_217__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4044) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2705 ( .A(
        mem_stage_inst_dmem_ram_217__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4045) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2704 ( .A(
        mem_stage_inst_dmem_ram_217__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4046) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2703 ( .A(
        mem_stage_inst_dmem_ram_217__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4047) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2702 ( .A(
        mem_stage_inst_dmem_ram_217__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4048) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2701 ( .A(
        mem_stage_inst_dmem_ram_217__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4049) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2700 ( .A(
        mem_stage_inst_dmem_ram_217__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4050) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2699 ( .A(
        mem_stage_inst_dmem_ram_217__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4051) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2698 ( .A(
        mem_stage_inst_dmem_ram_217__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5758), .Y(mem_stage_inst_dmem_n4052) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2697 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5757) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2696 ( .A(
        mem_stage_inst_dmem_ram_218__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4053) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2695 ( .A(
        mem_stage_inst_dmem_ram_218__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4054) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2694 ( .A(
        mem_stage_inst_dmem_ram_218__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4055) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2693 ( .A(
        mem_stage_inst_dmem_ram_218__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4056) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2692 ( .A(
        mem_stage_inst_dmem_ram_218__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4057) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2691 ( .A(
        mem_stage_inst_dmem_ram_218__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4058) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2690 ( .A(
        mem_stage_inst_dmem_ram_218__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4059) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2689 ( .A(
        mem_stage_inst_dmem_ram_218__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4060) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2688 ( .A(
        mem_stage_inst_dmem_ram_218__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4061) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2687 ( .A(
        mem_stage_inst_dmem_ram_218__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4062) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2686 ( .A(
        mem_stage_inst_dmem_ram_218__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4063) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2685 ( .A(
        mem_stage_inst_dmem_ram_218__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4064) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2684 ( .A(
        mem_stage_inst_dmem_ram_218__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4065) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2683 ( .A(
        mem_stage_inst_dmem_ram_218__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4066) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2682 ( .A(
        mem_stage_inst_dmem_ram_218__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4067) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2681 ( .A(
        mem_stage_inst_dmem_ram_218__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5757), .Y(mem_stage_inst_dmem_n4068) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2680 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5756) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2679 ( .A(
        mem_stage_inst_dmem_ram_219__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4069) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2678 ( .A(
        mem_stage_inst_dmem_ram_219__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4070) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2677 ( .A(
        mem_stage_inst_dmem_ram_219__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4071) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2676 ( .A(
        mem_stage_inst_dmem_ram_219__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4072) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2675 ( .A(
        mem_stage_inst_dmem_ram_219__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4073) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2674 ( .A(
        mem_stage_inst_dmem_ram_219__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4074) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2673 ( .A(
        mem_stage_inst_dmem_ram_219__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4075) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2672 ( .A(
        mem_stage_inst_dmem_ram_219__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4076) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2671 ( .A(
        mem_stage_inst_dmem_ram_219__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4077) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2670 ( .A(
        mem_stage_inst_dmem_ram_219__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4078) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2669 ( .A(
        mem_stage_inst_dmem_ram_219__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4079) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2668 ( .A(
        mem_stage_inst_dmem_ram_219__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4080) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2667 ( .A(
        mem_stage_inst_dmem_ram_219__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4081) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2666 ( .A(
        mem_stage_inst_dmem_ram_219__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4082) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2665 ( .A(
        mem_stage_inst_dmem_ram_219__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4083) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2664 ( .A(
        mem_stage_inst_dmem_ram_219__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5756), .Y(mem_stage_inst_dmem_n4084) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2663 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5755) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2662 ( .A(
        mem_stage_inst_dmem_ram_220__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4085) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2661 ( .A(
        mem_stage_inst_dmem_ram_220__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4086) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2660 ( .A(
        mem_stage_inst_dmem_ram_220__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4087) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2659 ( .A(
        mem_stage_inst_dmem_ram_220__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4088) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2658 ( .A(
        mem_stage_inst_dmem_ram_220__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4089) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2657 ( .A(
        mem_stage_inst_dmem_ram_220__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4090) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2656 ( .A(
        mem_stage_inst_dmem_ram_220__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4091) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2655 ( .A(
        mem_stage_inst_dmem_ram_220__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4092) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2654 ( .A(
        mem_stage_inst_dmem_ram_220__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4093) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2653 ( .A(
        mem_stage_inst_dmem_ram_220__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4094) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2652 ( .A(
        mem_stage_inst_dmem_ram_220__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4095) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2651 ( .A(
        mem_stage_inst_dmem_ram_220__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4096) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2650 ( .A(
        mem_stage_inst_dmem_ram_220__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4097) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2649 ( .A(
        mem_stage_inst_dmem_ram_220__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4098) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2648 ( .A(
        mem_stage_inst_dmem_ram_220__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4099) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2647 ( .A(
        mem_stage_inst_dmem_ram_220__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5755), .Y(mem_stage_inst_dmem_n4100) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2646 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5754) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2645 ( .A(
        mem_stage_inst_dmem_ram_221__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4101) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2644 ( .A(
        mem_stage_inst_dmem_ram_221__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4102) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2643 ( .A(
        mem_stage_inst_dmem_ram_221__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4103) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2642 ( .A(
        mem_stage_inst_dmem_ram_221__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4104) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2641 ( .A(
        mem_stage_inst_dmem_ram_221__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4105) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2640 ( .A(
        mem_stage_inst_dmem_ram_221__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4106) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2639 ( .A(
        mem_stage_inst_dmem_ram_221__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4107) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2638 ( .A(
        mem_stage_inst_dmem_ram_221__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4108) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2637 ( .A(
        mem_stage_inst_dmem_ram_221__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4109) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2636 ( .A(
        mem_stage_inst_dmem_ram_221__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4110) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2635 ( .A(
        mem_stage_inst_dmem_ram_221__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4111) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2634 ( .A(
        mem_stage_inst_dmem_ram_221__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4112) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2633 ( .A(
        mem_stage_inst_dmem_ram_221__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4113) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2632 ( .A(
        mem_stage_inst_dmem_ram_221__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4114) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2631 ( .A(
        mem_stage_inst_dmem_ram_221__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4115) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2630 ( .A(
        mem_stage_inst_dmem_ram_221__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5754), .Y(mem_stage_inst_dmem_n4116) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2629 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5753) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2628 ( .A(
        mem_stage_inst_dmem_ram_222__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4117) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2627 ( .A(
        mem_stage_inst_dmem_ram_222__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4118) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2626 ( .A(
        mem_stage_inst_dmem_ram_222__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4119) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2625 ( .A(
        mem_stage_inst_dmem_ram_222__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4120) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2624 ( .A(
        mem_stage_inst_dmem_ram_222__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4121) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2623 ( .A(
        mem_stage_inst_dmem_ram_222__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4122) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2622 ( .A(
        mem_stage_inst_dmem_ram_222__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4123) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2621 ( .A(
        mem_stage_inst_dmem_ram_222__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4124) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2620 ( .A(
        mem_stage_inst_dmem_ram_222__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4125) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2619 ( .A(
        mem_stage_inst_dmem_ram_222__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4126) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2618 ( .A(
        mem_stage_inst_dmem_ram_222__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4127) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2617 ( .A(
        mem_stage_inst_dmem_ram_222__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4128) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2616 ( .A(
        mem_stage_inst_dmem_ram_222__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4129) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2615 ( .A(
        mem_stage_inst_dmem_ram_222__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4130) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2614 ( .A(
        mem_stage_inst_dmem_ram_222__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4131) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2613 ( .A(
        mem_stage_inst_dmem_ram_222__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5753), .Y(mem_stage_inst_dmem_n4132) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2612 ( .A(mem_stage_inst_dmem_n5752), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5751) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2611 ( .A(
        mem_stage_inst_dmem_ram_223__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4133) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2610 ( .A(
        mem_stage_inst_dmem_ram_223__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4134) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2609 ( .A(
        mem_stage_inst_dmem_ram_223__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4135) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2608 ( .A(
        mem_stage_inst_dmem_ram_223__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4136) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2607 ( .A(
        mem_stage_inst_dmem_ram_223__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4137) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2606 ( .A(
        mem_stage_inst_dmem_ram_223__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4138) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2605 ( .A(
        mem_stage_inst_dmem_ram_223__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4139) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2604 ( .A(
        mem_stage_inst_dmem_ram_223__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4140) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2603 ( .A(
        mem_stage_inst_dmem_ram_223__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4141) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2602 ( .A(
        mem_stage_inst_dmem_ram_223__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4142) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2601 ( .A(
        mem_stage_inst_dmem_ram_223__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4143) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2600 ( .A(
        mem_stage_inst_dmem_ram_223__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4144) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2599 ( .A(
        mem_stage_inst_dmem_ram_223__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4145) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2598 ( .A(
        mem_stage_inst_dmem_ram_223__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4146) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2597 ( .A(
        mem_stage_inst_dmem_ram_223__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4147) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2596 ( .A(
        mem_stage_inst_dmem_ram_223__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5751), .Y(mem_stage_inst_dmem_n4148) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2595 ( .A(mem_stage_inst_dmem_n5750), 
        .B(mem_stage_inst_dmem_n5731), .Y(mem_stage_inst_dmem_n5734) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2594 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5749) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2593 ( .A(
        mem_stage_inst_dmem_ram_224__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4149) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2592 ( .A(
        mem_stage_inst_dmem_ram_224__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4150) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2591 ( .A(
        mem_stage_inst_dmem_ram_224__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4151) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2590 ( .A(
        mem_stage_inst_dmem_ram_224__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4152) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2589 ( .A(
        mem_stage_inst_dmem_ram_224__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4153) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2588 ( .A(
        mem_stage_inst_dmem_ram_224__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4154) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2587 ( .A(
        mem_stage_inst_dmem_ram_224__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4155) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2586 ( .A(
        mem_stage_inst_dmem_ram_224__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4156) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2585 ( .A(
        mem_stage_inst_dmem_ram_224__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4157) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2584 ( .A(
        mem_stage_inst_dmem_ram_224__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4158) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2583 ( .A(
        mem_stage_inst_dmem_ram_224__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4159) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2582 ( .A(
        mem_stage_inst_dmem_ram_224__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4160) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2581 ( .A(
        mem_stage_inst_dmem_ram_224__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4161) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2580 ( .A(
        mem_stage_inst_dmem_ram_224__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4162) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2579 ( .A(
        mem_stage_inst_dmem_ram_224__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4163) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2578 ( .A(
        mem_stage_inst_dmem_ram_224__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5749), .Y(mem_stage_inst_dmem_n4164) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2577 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5748) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2576 ( .A(
        mem_stage_inst_dmem_ram_225__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4165) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2575 ( .A(
        mem_stage_inst_dmem_ram_225__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4166) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2574 ( .A(
        mem_stage_inst_dmem_ram_225__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4167) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2573 ( .A(
        mem_stage_inst_dmem_ram_225__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4168) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2572 ( .A(
        mem_stage_inst_dmem_ram_225__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4169) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2571 ( .A(
        mem_stage_inst_dmem_ram_225__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4170) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2570 ( .A(
        mem_stage_inst_dmem_ram_225__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4171) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2569 ( .A(
        mem_stage_inst_dmem_ram_225__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4172) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2568 ( .A(
        mem_stage_inst_dmem_ram_225__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4173) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2567 ( .A(
        mem_stage_inst_dmem_ram_225__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4174) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2566 ( .A(
        mem_stage_inst_dmem_ram_225__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4175) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2565 ( .A(
        mem_stage_inst_dmem_ram_225__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4176) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2564 ( .A(
        mem_stage_inst_dmem_ram_225__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4177) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2563 ( .A(
        mem_stage_inst_dmem_ram_225__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4178) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2562 ( .A(
        mem_stage_inst_dmem_ram_225__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4179) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2561 ( .A(
        mem_stage_inst_dmem_ram_225__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5748), .Y(mem_stage_inst_dmem_n4180) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2560 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5747) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2559 ( .A(
        mem_stage_inst_dmem_ram_226__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4181) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2558 ( .A(
        mem_stage_inst_dmem_ram_226__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4182) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2557 ( .A(
        mem_stage_inst_dmem_ram_226__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4183) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2556 ( .A(
        mem_stage_inst_dmem_ram_226__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4184) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2555 ( .A(
        mem_stage_inst_dmem_ram_226__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4185) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2554 ( .A(
        mem_stage_inst_dmem_ram_226__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4186) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2553 ( .A(
        mem_stage_inst_dmem_ram_226__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4187) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2552 ( .A(
        mem_stage_inst_dmem_ram_226__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4188) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2551 ( .A(
        mem_stage_inst_dmem_ram_226__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4189) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2550 ( .A(
        mem_stage_inst_dmem_ram_226__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4190) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2549 ( .A(
        mem_stage_inst_dmem_ram_226__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4191) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2548 ( .A(
        mem_stage_inst_dmem_ram_226__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4192) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2547 ( .A(
        mem_stage_inst_dmem_ram_226__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4193) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2546 ( .A(
        mem_stage_inst_dmem_ram_226__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4194) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2545 ( .A(
        mem_stage_inst_dmem_ram_226__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4195) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2544 ( .A(
        mem_stage_inst_dmem_ram_226__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5747), .Y(mem_stage_inst_dmem_n4196) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2543 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5746) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2542 ( .A(
        mem_stage_inst_dmem_ram_227__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4197) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2541 ( .A(
        mem_stage_inst_dmem_ram_227__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4198) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2540 ( .A(
        mem_stage_inst_dmem_ram_227__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4199) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2539 ( .A(
        mem_stage_inst_dmem_ram_227__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4200) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2538 ( .A(
        mem_stage_inst_dmem_ram_227__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4201) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2537 ( .A(
        mem_stage_inst_dmem_ram_227__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4202) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2536 ( .A(
        mem_stage_inst_dmem_ram_227__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4203) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2535 ( .A(
        mem_stage_inst_dmem_ram_227__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4204) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2534 ( .A(
        mem_stage_inst_dmem_ram_227__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4205) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2533 ( .A(
        mem_stage_inst_dmem_ram_227__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4206) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2532 ( .A(
        mem_stage_inst_dmem_ram_227__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4207) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2531 ( .A(
        mem_stage_inst_dmem_ram_227__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4208) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2530 ( .A(
        mem_stage_inst_dmem_ram_227__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4209) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2529 ( .A(
        mem_stage_inst_dmem_ram_227__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4210) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2528 ( .A(
        mem_stage_inst_dmem_ram_227__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4211) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2527 ( .A(
        mem_stage_inst_dmem_ram_227__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5746), .Y(mem_stage_inst_dmem_n4212) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2526 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5745) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2525 ( .A(
        mem_stage_inst_dmem_ram_228__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4213) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2524 ( .A(
        mem_stage_inst_dmem_ram_228__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4214) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2523 ( .A(
        mem_stage_inst_dmem_ram_228__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4215) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2522 ( .A(
        mem_stage_inst_dmem_ram_228__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4216) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2521 ( .A(
        mem_stage_inst_dmem_ram_228__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4217) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2520 ( .A(
        mem_stage_inst_dmem_ram_228__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4218) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2519 ( .A(
        mem_stage_inst_dmem_ram_228__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4219) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2518 ( .A(
        mem_stage_inst_dmem_ram_228__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4220) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2517 ( .A(
        mem_stage_inst_dmem_ram_228__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4221) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2516 ( .A(
        mem_stage_inst_dmem_ram_228__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4222) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2515 ( .A(
        mem_stage_inst_dmem_ram_228__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4223) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2514 ( .A(
        mem_stage_inst_dmem_ram_228__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4224) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2513 ( .A(
        mem_stage_inst_dmem_ram_228__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4225) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2512 ( .A(
        mem_stage_inst_dmem_ram_228__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4226) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2511 ( .A(
        mem_stage_inst_dmem_ram_228__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4227) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2510 ( .A(
        mem_stage_inst_dmem_ram_228__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5745), .Y(mem_stage_inst_dmem_n4228) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2509 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5744) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2508 ( .A(
        mem_stage_inst_dmem_ram_229__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4229) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2507 ( .A(
        mem_stage_inst_dmem_ram_229__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4230) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2506 ( .A(
        mem_stage_inst_dmem_ram_229__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4231) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2505 ( .A(
        mem_stage_inst_dmem_ram_229__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4232) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2504 ( .A(
        mem_stage_inst_dmem_ram_229__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4233) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2503 ( .A(
        mem_stage_inst_dmem_ram_229__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4234) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2502 ( .A(
        mem_stage_inst_dmem_ram_229__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4235) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2501 ( .A(
        mem_stage_inst_dmem_ram_229__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4236) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2500 ( .A(
        mem_stage_inst_dmem_ram_229__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4237) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2499 ( .A(
        mem_stage_inst_dmem_ram_229__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4238) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2498 ( .A(
        mem_stage_inst_dmem_ram_229__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4239) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2497 ( .A(
        mem_stage_inst_dmem_ram_229__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4240) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2496 ( .A(
        mem_stage_inst_dmem_ram_229__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4241) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2495 ( .A(
        mem_stage_inst_dmem_ram_229__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4242) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2494 ( .A(
        mem_stage_inst_dmem_ram_229__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4243) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2493 ( .A(
        mem_stage_inst_dmem_ram_229__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5744), .Y(mem_stage_inst_dmem_n4244) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2492 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5743) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2491 ( .A(
        mem_stage_inst_dmem_ram_230__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4245) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2490 ( .A(
        mem_stage_inst_dmem_ram_230__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4246) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2489 ( .A(
        mem_stage_inst_dmem_ram_230__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4247) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2488 ( .A(
        mem_stage_inst_dmem_ram_230__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4248) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2487 ( .A(
        mem_stage_inst_dmem_ram_230__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4249) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2486 ( .A(
        mem_stage_inst_dmem_ram_230__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4250) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2485 ( .A(
        mem_stage_inst_dmem_ram_230__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4251) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2484 ( .A(
        mem_stage_inst_dmem_ram_230__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4252) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2483 ( .A(
        mem_stage_inst_dmem_ram_230__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4253) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2482 ( .A(
        mem_stage_inst_dmem_ram_230__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4254) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2481 ( .A(
        mem_stage_inst_dmem_ram_230__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4255) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2480 ( .A(
        mem_stage_inst_dmem_ram_230__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4256) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2479 ( .A(
        mem_stage_inst_dmem_ram_230__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4257) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2478 ( .A(
        mem_stage_inst_dmem_ram_230__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4258) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2477 ( .A(
        mem_stage_inst_dmem_ram_230__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4259) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2476 ( .A(
        mem_stage_inst_dmem_ram_230__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5743), .Y(mem_stage_inst_dmem_n4260) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2475 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5742) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2474 ( .A(
        mem_stage_inst_dmem_ram_231__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4261) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2473 ( .A(
        mem_stage_inst_dmem_ram_231__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4262) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2472 ( .A(
        mem_stage_inst_dmem_ram_231__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4263) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2471 ( .A(
        mem_stage_inst_dmem_ram_231__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4264) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2470 ( .A(
        mem_stage_inst_dmem_ram_231__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4265) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2469 ( .A(
        mem_stage_inst_dmem_ram_231__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4266) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2468 ( .A(
        mem_stage_inst_dmem_ram_231__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4267) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2467 ( .A(
        mem_stage_inst_dmem_ram_231__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4268) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2466 ( .A(
        mem_stage_inst_dmem_ram_231__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4269) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2465 ( .A(
        mem_stage_inst_dmem_ram_231__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4270) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2464 ( .A(
        mem_stage_inst_dmem_ram_231__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4271) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2463 ( .A(
        mem_stage_inst_dmem_ram_231__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4272) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2462 ( .A(
        mem_stage_inst_dmem_ram_231__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4273) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2461 ( .A(
        mem_stage_inst_dmem_ram_231__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4274) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2460 ( .A(
        mem_stage_inst_dmem_ram_231__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4275) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2459 ( .A(
        mem_stage_inst_dmem_ram_231__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5742), .Y(mem_stage_inst_dmem_n4276) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2458 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5741) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2457 ( .A(
        mem_stage_inst_dmem_ram_232__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4277) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2456 ( .A(
        mem_stage_inst_dmem_ram_232__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4278) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2455 ( .A(
        mem_stage_inst_dmem_ram_232__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4279) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2454 ( .A(
        mem_stage_inst_dmem_ram_232__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4280) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2453 ( .A(
        mem_stage_inst_dmem_ram_232__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4281) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2452 ( .A(
        mem_stage_inst_dmem_ram_232__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4282) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2451 ( .A(
        mem_stage_inst_dmem_ram_232__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4283) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2450 ( .A(
        mem_stage_inst_dmem_ram_232__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4284) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2449 ( .A(
        mem_stage_inst_dmem_ram_232__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4285) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2448 ( .A(
        mem_stage_inst_dmem_ram_232__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4286) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2447 ( .A(
        mem_stage_inst_dmem_ram_232__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4287) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2446 ( .A(
        mem_stage_inst_dmem_ram_232__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4288) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2445 ( .A(
        mem_stage_inst_dmem_ram_232__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4289) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2444 ( .A(
        mem_stage_inst_dmem_ram_232__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4290) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2443 ( .A(
        mem_stage_inst_dmem_ram_232__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4291) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2442 ( .A(
        mem_stage_inst_dmem_ram_232__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5741), .Y(mem_stage_inst_dmem_n4292) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2441 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5740) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2440 ( .A(
        mem_stage_inst_dmem_ram_233__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4293) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2439 ( .A(
        mem_stage_inst_dmem_ram_233__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4294) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2438 ( .A(
        mem_stage_inst_dmem_ram_233__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4295) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2437 ( .A(
        mem_stage_inst_dmem_ram_233__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4296) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2436 ( .A(
        mem_stage_inst_dmem_ram_233__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4297) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2435 ( .A(
        mem_stage_inst_dmem_ram_233__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4298) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2434 ( .A(
        mem_stage_inst_dmem_ram_233__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4299) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2433 ( .A(
        mem_stage_inst_dmem_ram_233__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4300) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2432 ( .A(
        mem_stage_inst_dmem_ram_233__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4301) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2431 ( .A(
        mem_stage_inst_dmem_ram_233__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4302) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2430 ( .A(
        mem_stage_inst_dmem_ram_233__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4303) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2429 ( .A(
        mem_stage_inst_dmem_ram_233__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4304) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2428 ( .A(
        mem_stage_inst_dmem_ram_233__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4305) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2427 ( .A(
        mem_stage_inst_dmem_ram_233__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4306) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2426 ( .A(
        mem_stage_inst_dmem_ram_233__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4307) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2425 ( .A(
        mem_stage_inst_dmem_ram_233__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5740), .Y(mem_stage_inst_dmem_n4308) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2424 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5739) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2423 ( .A(
        mem_stage_inst_dmem_ram_234__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4309) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2422 ( .A(
        mem_stage_inst_dmem_ram_234__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4310) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2421 ( .A(
        mem_stage_inst_dmem_ram_234__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4311) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2420 ( .A(
        mem_stage_inst_dmem_ram_234__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4312) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2419 ( .A(
        mem_stage_inst_dmem_ram_234__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4313) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2418 ( .A(
        mem_stage_inst_dmem_ram_234__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4314) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2417 ( .A(
        mem_stage_inst_dmem_ram_234__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4315) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2416 ( .A(
        mem_stage_inst_dmem_ram_234__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4316) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2415 ( .A(
        mem_stage_inst_dmem_ram_234__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4317) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2414 ( .A(
        mem_stage_inst_dmem_ram_234__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4318) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2413 ( .A(
        mem_stage_inst_dmem_ram_234__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4319) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2412 ( .A(
        mem_stage_inst_dmem_ram_234__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4320) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2411 ( .A(
        mem_stage_inst_dmem_ram_234__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4321) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2410 ( .A(
        mem_stage_inst_dmem_ram_234__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4322) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2409 ( .A(
        mem_stage_inst_dmem_ram_234__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4323) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2408 ( .A(
        mem_stage_inst_dmem_ram_234__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5739), .Y(mem_stage_inst_dmem_n4324) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2407 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5738) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2406 ( .A(
        mem_stage_inst_dmem_ram_235__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4325) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2405 ( .A(
        mem_stage_inst_dmem_ram_235__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4326) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2404 ( .A(
        mem_stage_inst_dmem_ram_235__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4327) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2403 ( .A(
        mem_stage_inst_dmem_ram_235__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4328) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2402 ( .A(
        mem_stage_inst_dmem_ram_235__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4329) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2401 ( .A(
        mem_stage_inst_dmem_ram_235__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4330) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2400 ( .A(
        mem_stage_inst_dmem_ram_235__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4331) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2399 ( .A(
        mem_stage_inst_dmem_ram_235__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4332) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2398 ( .A(
        mem_stage_inst_dmem_ram_235__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4333) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2397 ( .A(
        mem_stage_inst_dmem_ram_235__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4334) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2396 ( .A(
        mem_stage_inst_dmem_ram_235__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4335) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2395 ( .A(
        mem_stage_inst_dmem_ram_235__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4336) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2394 ( .A(
        mem_stage_inst_dmem_ram_235__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4337) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2393 ( .A(
        mem_stage_inst_dmem_ram_235__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4338) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2392 ( .A(
        mem_stage_inst_dmem_ram_235__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4339) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2391 ( .A(
        mem_stage_inst_dmem_ram_235__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5738), .Y(mem_stage_inst_dmem_n4340) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2390 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5737) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2389 ( .A(
        mem_stage_inst_dmem_ram_236__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4341) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2388 ( .A(
        mem_stage_inst_dmem_ram_236__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4342) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2387 ( .A(
        mem_stage_inst_dmem_ram_236__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4343) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2386 ( .A(
        mem_stage_inst_dmem_ram_236__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4344) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2385 ( .A(
        mem_stage_inst_dmem_ram_236__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4345) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2384 ( .A(
        mem_stage_inst_dmem_ram_236__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4346) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2383 ( .A(
        mem_stage_inst_dmem_ram_236__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4347) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2382 ( .A(
        mem_stage_inst_dmem_ram_236__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4348) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2381 ( .A(
        mem_stage_inst_dmem_ram_236__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4349) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2380 ( .A(
        mem_stage_inst_dmem_ram_236__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4350) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2379 ( .A(
        mem_stage_inst_dmem_ram_236__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4351) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2378 ( .A(
        mem_stage_inst_dmem_ram_236__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4352) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2377 ( .A(
        mem_stage_inst_dmem_ram_236__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4353) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2376 ( .A(
        mem_stage_inst_dmem_ram_236__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4354) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2375 ( .A(
        mem_stage_inst_dmem_ram_236__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4355) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2374 ( .A(
        mem_stage_inst_dmem_ram_236__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5737), .Y(mem_stage_inst_dmem_n4356) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2373 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5736) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2372 ( .A(
        mem_stage_inst_dmem_ram_237__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4357) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2371 ( .A(
        mem_stage_inst_dmem_ram_237__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4358) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2370 ( .A(
        mem_stage_inst_dmem_ram_237__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4359) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2369 ( .A(
        mem_stage_inst_dmem_ram_237__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4360) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2368 ( .A(
        mem_stage_inst_dmem_ram_237__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4361) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2367 ( .A(
        mem_stage_inst_dmem_ram_237__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4362) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2366 ( .A(
        mem_stage_inst_dmem_ram_237__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4363) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2365 ( .A(
        mem_stage_inst_dmem_ram_237__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4364) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2364 ( .A(
        mem_stage_inst_dmem_ram_237__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4365) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2363 ( .A(
        mem_stage_inst_dmem_ram_237__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4366) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2362 ( .A(
        mem_stage_inst_dmem_ram_237__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4367) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2361 ( .A(
        mem_stage_inst_dmem_ram_237__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4368) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2360 ( .A(
        mem_stage_inst_dmem_ram_237__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4369) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2359 ( .A(
        mem_stage_inst_dmem_ram_237__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4370) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2358 ( .A(
        mem_stage_inst_dmem_ram_237__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4371) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2357 ( .A(
        mem_stage_inst_dmem_ram_237__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5736), .Y(mem_stage_inst_dmem_n4372) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2356 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5735) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2355 ( .A(
        mem_stage_inst_dmem_ram_238__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4373) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2354 ( .A(
        mem_stage_inst_dmem_ram_238__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4374) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2353 ( .A(
        mem_stage_inst_dmem_ram_238__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4375) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2352 ( .A(
        mem_stage_inst_dmem_ram_238__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4376) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2351 ( .A(
        mem_stage_inst_dmem_ram_238__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4377) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2350 ( .A(
        mem_stage_inst_dmem_ram_238__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4378) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2349 ( .A(
        mem_stage_inst_dmem_ram_238__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4379) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2348 ( .A(
        mem_stage_inst_dmem_ram_238__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4380) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2347 ( .A(
        mem_stage_inst_dmem_ram_238__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4381) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2346 ( .A(
        mem_stage_inst_dmem_ram_238__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4382) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2345 ( .A(
        mem_stage_inst_dmem_ram_238__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4383) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2344 ( .A(
        mem_stage_inst_dmem_ram_238__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4384) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2343 ( .A(
        mem_stage_inst_dmem_ram_238__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4385) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2342 ( .A(
        mem_stage_inst_dmem_ram_238__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4386) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2341 ( .A(
        mem_stage_inst_dmem_ram_238__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4387) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2340 ( .A(
        mem_stage_inst_dmem_ram_238__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5735), .Y(mem_stage_inst_dmem_n4388) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2339 ( .A(mem_stage_inst_dmem_n5734), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5733) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2338 ( .A(
        mem_stage_inst_dmem_ram_239__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4389) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2337 ( .A(
        mem_stage_inst_dmem_ram_239__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4390) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2336 ( .A(
        mem_stage_inst_dmem_ram_239__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4391) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2335 ( .A(
        mem_stage_inst_dmem_ram_239__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4392) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2334 ( .A(
        mem_stage_inst_dmem_ram_239__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4393) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2333 ( .A(
        mem_stage_inst_dmem_ram_239__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4394) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2332 ( .A(
        mem_stage_inst_dmem_ram_239__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4395) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2331 ( .A(
        mem_stage_inst_dmem_ram_239__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4396) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2330 ( .A(
        mem_stage_inst_dmem_ram_239__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4397) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2329 ( .A(
        mem_stage_inst_dmem_ram_239__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4398) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2328 ( .A(
        mem_stage_inst_dmem_ram_239__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4399) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2327 ( .A(
        mem_stage_inst_dmem_ram_239__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4400) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2326 ( .A(
        mem_stage_inst_dmem_ram_239__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4401) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2325 ( .A(
        mem_stage_inst_dmem_ram_239__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4402) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2324 ( .A(
        mem_stage_inst_dmem_ram_239__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4403) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2323 ( .A(
        mem_stage_inst_dmem_ram_239__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5733), .Y(mem_stage_inst_dmem_n4404) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2322 ( .A(mem_stage_inst_dmem_n5731), 
        .B(mem_stage_inst_dmem_n5732), .Y(mem_stage_inst_dmem_n5715) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2321 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5730) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2320 ( .A(
        mem_stage_inst_dmem_ram_240__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4405) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2319 ( .A(
        mem_stage_inst_dmem_ram_240__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4406) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2318 ( .A(
        mem_stage_inst_dmem_ram_240__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4407) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2317 ( .A(
        mem_stage_inst_dmem_ram_240__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4408) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2316 ( .A(
        mem_stage_inst_dmem_ram_240__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4409) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2315 ( .A(
        mem_stage_inst_dmem_ram_240__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4410) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2314 ( .A(
        mem_stage_inst_dmem_ram_240__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4411) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2313 ( .A(
        mem_stage_inst_dmem_ram_240__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4412) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2312 ( .A(
        mem_stage_inst_dmem_ram_240__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4413) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2311 ( .A(
        mem_stage_inst_dmem_ram_240__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4414) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2310 ( .A(
        mem_stage_inst_dmem_ram_240__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4415) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2309 ( .A(
        mem_stage_inst_dmem_ram_240__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4416) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2308 ( .A(
        mem_stage_inst_dmem_ram_240__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4417) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2307 ( .A(
        mem_stage_inst_dmem_ram_240__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4418) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2306 ( .A(
        mem_stage_inst_dmem_ram_240__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4419) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2305 ( .A(
        mem_stage_inst_dmem_ram_240__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5730), .Y(mem_stage_inst_dmem_n4420) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2304 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5729) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2303 ( .A(
        mem_stage_inst_dmem_ram_241__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4421) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2302 ( .A(
        mem_stage_inst_dmem_ram_241__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4422) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2301 ( .A(
        mem_stage_inst_dmem_ram_241__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4423) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2300 ( .A(
        mem_stage_inst_dmem_ram_241__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4424) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2299 ( .A(
        mem_stage_inst_dmem_ram_241__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4425) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2298 ( .A(
        mem_stage_inst_dmem_ram_241__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4426) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2297 ( .A(
        mem_stage_inst_dmem_ram_241__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4427) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2296 ( .A(
        mem_stage_inst_dmem_ram_241__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4428) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2295 ( .A(
        mem_stage_inst_dmem_ram_241__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4429) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2294 ( .A(
        mem_stage_inst_dmem_ram_241__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4430) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2293 ( .A(
        mem_stage_inst_dmem_ram_241__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4431) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2292 ( .A(
        mem_stage_inst_dmem_ram_241__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4432) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2291 ( .A(
        mem_stage_inst_dmem_ram_241__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4433) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2290 ( .A(
        mem_stage_inst_dmem_ram_241__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4434) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2289 ( .A(
        mem_stage_inst_dmem_ram_241__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4435) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2288 ( .A(
        mem_stage_inst_dmem_ram_241__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5729), .Y(mem_stage_inst_dmem_n4436) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2287 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5728) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2286 ( .A(
        mem_stage_inst_dmem_ram_242__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4437) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2285 ( .A(
        mem_stage_inst_dmem_ram_242__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4438) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2284 ( .A(
        mem_stage_inst_dmem_ram_242__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4439) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2283 ( .A(
        mem_stage_inst_dmem_ram_242__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4440) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2282 ( .A(
        mem_stage_inst_dmem_ram_242__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4441) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2281 ( .A(
        mem_stage_inst_dmem_ram_242__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4442) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2280 ( .A(
        mem_stage_inst_dmem_ram_242__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4443) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2279 ( .A(
        mem_stage_inst_dmem_ram_242__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4444) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2278 ( .A(
        mem_stage_inst_dmem_ram_242__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4445) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2277 ( .A(
        mem_stage_inst_dmem_ram_242__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4446) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2276 ( .A(
        mem_stage_inst_dmem_ram_242__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4447) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2275 ( .A(
        mem_stage_inst_dmem_ram_242__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4448) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2274 ( .A(
        mem_stage_inst_dmem_ram_242__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4449) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2273 ( .A(
        mem_stage_inst_dmem_ram_242__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4450) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2272 ( .A(
        mem_stage_inst_dmem_ram_242__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4451) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2271 ( .A(
        mem_stage_inst_dmem_ram_242__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5728), .Y(mem_stage_inst_dmem_n4452) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2270 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5727) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2269 ( .A(
        mem_stage_inst_dmem_ram_243__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4453) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2268 ( .A(
        mem_stage_inst_dmem_ram_243__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4454) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2267 ( .A(
        mem_stage_inst_dmem_ram_243__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4455) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2266 ( .A(
        mem_stage_inst_dmem_ram_243__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4456) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2265 ( .A(
        mem_stage_inst_dmem_ram_243__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4457) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2264 ( .A(
        mem_stage_inst_dmem_ram_243__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4458) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2263 ( .A(
        mem_stage_inst_dmem_ram_243__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4459) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2262 ( .A(
        mem_stage_inst_dmem_ram_243__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4460) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2261 ( .A(
        mem_stage_inst_dmem_ram_243__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4461) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2260 ( .A(
        mem_stage_inst_dmem_ram_243__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4462) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2259 ( .A(
        mem_stage_inst_dmem_ram_243__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4463) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2258 ( .A(
        mem_stage_inst_dmem_ram_243__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4464) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2257 ( .A(
        mem_stage_inst_dmem_ram_243__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4465) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2256 ( .A(
        mem_stage_inst_dmem_ram_243__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4466) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2255 ( .A(
        mem_stage_inst_dmem_ram_243__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4467) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2254 ( .A(
        mem_stage_inst_dmem_ram_243__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5727), .Y(mem_stage_inst_dmem_n4468) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2253 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5726) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2252 ( .A(
        mem_stage_inst_dmem_ram_244__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4469) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2251 ( .A(
        mem_stage_inst_dmem_ram_244__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4470) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2250 ( .A(
        mem_stage_inst_dmem_ram_244__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4471) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2249 ( .A(
        mem_stage_inst_dmem_ram_244__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4472) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2248 ( .A(
        mem_stage_inst_dmem_ram_244__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4473) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2247 ( .A(
        mem_stage_inst_dmem_ram_244__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4474) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2246 ( .A(
        mem_stage_inst_dmem_ram_244__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4475) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2245 ( .A(
        mem_stage_inst_dmem_ram_244__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4476) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2244 ( .A(
        mem_stage_inst_dmem_ram_244__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4477) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2243 ( .A(
        mem_stage_inst_dmem_ram_244__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4478) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2242 ( .A(
        mem_stage_inst_dmem_ram_244__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4479) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2241 ( .A(
        mem_stage_inst_dmem_ram_244__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4480) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2240 ( .A(
        mem_stage_inst_dmem_ram_244__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4481) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2239 ( .A(
        mem_stage_inst_dmem_ram_244__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4482) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2238 ( .A(
        mem_stage_inst_dmem_ram_244__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4483) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2237 ( .A(
        mem_stage_inst_dmem_ram_244__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5726), .Y(mem_stage_inst_dmem_n4484) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2236 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5725) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2235 ( .A(
        mem_stage_inst_dmem_ram_245__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4485) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2234 ( .A(
        mem_stage_inst_dmem_ram_245__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4486) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2233 ( .A(
        mem_stage_inst_dmem_ram_245__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4487) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2232 ( .A(
        mem_stage_inst_dmem_ram_245__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4488) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2231 ( .A(
        mem_stage_inst_dmem_ram_245__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4489) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2230 ( .A(
        mem_stage_inst_dmem_ram_245__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4490) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2229 ( .A(
        mem_stage_inst_dmem_ram_245__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4491) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2228 ( .A(
        mem_stage_inst_dmem_ram_245__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4492) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2227 ( .A(
        mem_stage_inst_dmem_ram_245__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4493) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2226 ( .A(
        mem_stage_inst_dmem_ram_245__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4494) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2225 ( .A(
        mem_stage_inst_dmem_ram_245__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4495) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2224 ( .A(
        mem_stage_inst_dmem_ram_245__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4496) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2223 ( .A(
        mem_stage_inst_dmem_ram_245__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4497) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2222 ( .A(
        mem_stage_inst_dmem_ram_245__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4498) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2221 ( .A(
        mem_stage_inst_dmem_ram_245__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4499) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2220 ( .A(
        mem_stage_inst_dmem_ram_245__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5725), .Y(mem_stage_inst_dmem_n4500) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2219 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5724) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2218 ( .A(
        mem_stage_inst_dmem_ram_246__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4501) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2217 ( .A(
        mem_stage_inst_dmem_ram_246__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4502) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2216 ( .A(
        mem_stage_inst_dmem_ram_246__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4503) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2215 ( .A(
        mem_stage_inst_dmem_ram_246__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4504) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2214 ( .A(
        mem_stage_inst_dmem_ram_246__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4505) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2213 ( .A(
        mem_stage_inst_dmem_ram_246__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4506) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2212 ( .A(
        mem_stage_inst_dmem_ram_246__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4507) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2211 ( .A(
        mem_stage_inst_dmem_ram_246__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4508) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2210 ( .A(
        mem_stage_inst_dmem_ram_246__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4509) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2209 ( .A(
        mem_stage_inst_dmem_ram_246__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4510) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2208 ( .A(
        mem_stage_inst_dmem_ram_246__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4511) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2207 ( .A(
        mem_stage_inst_dmem_ram_246__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4512) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2206 ( .A(
        mem_stage_inst_dmem_ram_246__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4513) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2205 ( .A(
        mem_stage_inst_dmem_ram_246__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4514) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2204 ( .A(
        mem_stage_inst_dmem_ram_246__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4515) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2203 ( .A(
        mem_stage_inst_dmem_ram_246__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5724), .Y(mem_stage_inst_dmem_n4516) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2202 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5723) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2201 ( .A(
        mem_stage_inst_dmem_ram_247__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4517) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2200 ( .A(
        mem_stage_inst_dmem_ram_247__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4518) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2199 ( .A(
        mem_stage_inst_dmem_ram_247__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4519) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2198 ( .A(
        mem_stage_inst_dmem_ram_247__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4520) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2197 ( .A(
        mem_stage_inst_dmem_ram_247__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4521) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2196 ( .A(
        mem_stage_inst_dmem_ram_247__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4522) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2195 ( .A(
        mem_stage_inst_dmem_ram_247__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4523) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2194 ( .A(
        mem_stage_inst_dmem_ram_247__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4524) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2193 ( .A(
        mem_stage_inst_dmem_ram_247__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4525) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2192 ( .A(
        mem_stage_inst_dmem_ram_247__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4526) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2191 ( .A(
        mem_stage_inst_dmem_ram_247__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4527) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2190 ( .A(
        mem_stage_inst_dmem_ram_247__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4528) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2189 ( .A(
        mem_stage_inst_dmem_ram_247__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4529) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2188 ( .A(
        mem_stage_inst_dmem_ram_247__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4530) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2187 ( .A(
        mem_stage_inst_dmem_ram_247__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4531) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2186 ( .A(
        mem_stage_inst_dmem_ram_247__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5723), .Y(mem_stage_inst_dmem_n4532) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2185 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5722) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2184 ( .A(
        mem_stage_inst_dmem_ram_248__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4533) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2183 ( .A(
        mem_stage_inst_dmem_ram_248__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4534) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2182 ( .A(
        mem_stage_inst_dmem_ram_248__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4535) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2181 ( .A(
        mem_stage_inst_dmem_ram_248__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4536) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2180 ( .A(
        mem_stage_inst_dmem_ram_248__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4537) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2179 ( .A(
        mem_stage_inst_dmem_ram_248__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4538) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2178 ( .A(
        mem_stage_inst_dmem_ram_248__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4539) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2177 ( .A(
        mem_stage_inst_dmem_ram_248__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4540) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2176 ( .A(
        mem_stage_inst_dmem_ram_248__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4541) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2175 ( .A(
        mem_stage_inst_dmem_ram_248__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4542) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2174 ( .A(
        mem_stage_inst_dmem_ram_248__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4543) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2173 ( .A(
        mem_stage_inst_dmem_ram_248__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4544) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2172 ( .A(
        mem_stage_inst_dmem_ram_248__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4545) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2171 ( .A(
        mem_stage_inst_dmem_ram_248__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4546) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2170 ( .A(
        mem_stage_inst_dmem_ram_248__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4547) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2169 ( .A(
        mem_stage_inst_dmem_ram_248__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5722), .Y(mem_stage_inst_dmem_n4548) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2168 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5721) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2167 ( .A(
        mem_stage_inst_dmem_ram_249__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4549) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2166 ( .A(
        mem_stage_inst_dmem_ram_249__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4550) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2165 ( .A(
        mem_stage_inst_dmem_ram_249__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4551) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2164 ( .A(
        mem_stage_inst_dmem_ram_249__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4552) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2163 ( .A(
        mem_stage_inst_dmem_ram_249__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4553) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2162 ( .A(
        mem_stage_inst_dmem_ram_249__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4554) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2161 ( .A(
        mem_stage_inst_dmem_ram_249__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4555) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2160 ( .A(
        mem_stage_inst_dmem_ram_249__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4556) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2159 ( .A(
        mem_stage_inst_dmem_ram_249__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4557) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2158 ( .A(
        mem_stage_inst_dmem_ram_249__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4558) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2157 ( .A(
        mem_stage_inst_dmem_ram_249__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4559) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2156 ( .A(
        mem_stage_inst_dmem_ram_249__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4560) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2155 ( .A(
        mem_stage_inst_dmem_ram_249__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4561) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2154 ( .A(
        mem_stage_inst_dmem_ram_249__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4562) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2153 ( .A(
        mem_stage_inst_dmem_ram_249__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4563) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2152 ( .A(
        mem_stage_inst_dmem_ram_249__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5721), .Y(mem_stage_inst_dmem_n4564) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2151 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5720) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2150 ( .A(
        mem_stage_inst_dmem_ram_250__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4565) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2149 ( .A(
        mem_stage_inst_dmem_ram_250__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4566) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2148 ( .A(
        mem_stage_inst_dmem_ram_250__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4567) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2147 ( .A(
        mem_stage_inst_dmem_ram_250__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4568) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2146 ( .A(
        mem_stage_inst_dmem_ram_250__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4569) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2145 ( .A(
        mem_stage_inst_dmem_ram_250__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4570) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2144 ( .A(
        mem_stage_inst_dmem_ram_250__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4571) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2143 ( .A(
        mem_stage_inst_dmem_ram_250__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4572) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2142 ( .A(
        mem_stage_inst_dmem_ram_250__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4573) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2141 ( .A(
        mem_stage_inst_dmem_ram_250__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4574) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2140 ( .A(
        mem_stage_inst_dmem_ram_250__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4575) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2139 ( .A(
        mem_stage_inst_dmem_ram_250__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4576) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2138 ( .A(
        mem_stage_inst_dmem_ram_250__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4577) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2137 ( .A(
        mem_stage_inst_dmem_ram_250__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4578) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2136 ( .A(
        mem_stage_inst_dmem_ram_250__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4579) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2135 ( .A(
        mem_stage_inst_dmem_ram_250__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5720), .Y(mem_stage_inst_dmem_n4580) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2134 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5719) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2133 ( .A(
        mem_stage_inst_dmem_ram_251__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4581) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2132 ( .A(
        mem_stage_inst_dmem_ram_251__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4582) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2131 ( .A(
        mem_stage_inst_dmem_ram_251__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4583) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2130 ( .A(
        mem_stage_inst_dmem_ram_251__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4584) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2129 ( .A(
        mem_stage_inst_dmem_ram_251__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4585) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2128 ( .A(
        mem_stage_inst_dmem_ram_251__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4586) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2127 ( .A(
        mem_stage_inst_dmem_ram_251__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4587) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2126 ( .A(
        mem_stage_inst_dmem_ram_251__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4588) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2125 ( .A(
        mem_stage_inst_dmem_ram_251__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4589) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2124 ( .A(
        mem_stage_inst_dmem_ram_251__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4590) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2123 ( .A(
        mem_stage_inst_dmem_ram_251__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4591) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2122 ( .A(
        mem_stage_inst_dmem_ram_251__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4592) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2121 ( .A(
        mem_stage_inst_dmem_ram_251__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4593) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2120 ( .A(
        mem_stage_inst_dmem_ram_251__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4594) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2119 ( .A(
        mem_stage_inst_dmem_ram_251__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4595) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2118 ( .A(
        mem_stage_inst_dmem_ram_251__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5719), .Y(mem_stage_inst_dmem_n4596) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2117 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5698), .Y(mem_stage_inst_dmem_n5718) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2116 ( .A(
        mem_stage_inst_dmem_ram_252__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4597) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2115 ( .A(
        mem_stage_inst_dmem_ram_252__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4598) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2114 ( .A(
        mem_stage_inst_dmem_ram_252__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4599) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2113 ( .A(
        mem_stage_inst_dmem_ram_252__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4600) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2112 ( .A(
        mem_stage_inst_dmem_ram_252__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4601) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2111 ( .A(
        mem_stage_inst_dmem_ram_252__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4602) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2110 ( .A(
        mem_stage_inst_dmem_ram_252__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4603) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2109 ( .A(
        mem_stage_inst_dmem_ram_252__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4604) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2108 ( .A(
        mem_stage_inst_dmem_ram_252__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4605) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2107 ( .A(
        mem_stage_inst_dmem_ram_252__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4606) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2106 ( .A(
        mem_stage_inst_dmem_ram_252__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4607) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2105 ( .A(
        mem_stage_inst_dmem_ram_252__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4608) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2104 ( .A(
        mem_stage_inst_dmem_ram_252__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4609) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2103 ( .A(
        mem_stage_inst_dmem_ram_252__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4610) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2102 ( .A(
        mem_stage_inst_dmem_ram_252__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4611) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2101 ( .A(
        mem_stage_inst_dmem_ram_252__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5718), .Y(mem_stage_inst_dmem_n4612) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2100 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5696), .Y(mem_stage_inst_dmem_n5717) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2099 ( .A(
        mem_stage_inst_dmem_ram_253__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4613) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2098 ( .A(
        mem_stage_inst_dmem_ram_253__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4614) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2097 ( .A(
        mem_stage_inst_dmem_ram_253__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4615) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2096 ( .A(
        mem_stage_inst_dmem_ram_253__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4616) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2095 ( .A(
        mem_stage_inst_dmem_ram_253__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4617) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2094 ( .A(
        mem_stage_inst_dmem_ram_253__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4618) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2093 ( .A(
        mem_stage_inst_dmem_ram_253__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4619) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2092 ( .A(
        mem_stage_inst_dmem_ram_253__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4620) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2091 ( .A(
        mem_stage_inst_dmem_ram_253__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4621) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2090 ( .A(
        mem_stage_inst_dmem_ram_253__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4622) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2089 ( .A(
        mem_stage_inst_dmem_ram_253__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4623) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2088 ( .A(
        mem_stage_inst_dmem_ram_253__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4624) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2087 ( .A(
        mem_stage_inst_dmem_ram_253__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4625) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2086 ( .A(
        mem_stage_inst_dmem_ram_253__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4626) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2085 ( .A(
        mem_stage_inst_dmem_ram_253__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4627) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2084 ( .A(
        mem_stage_inst_dmem_ram_253__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5717), .Y(mem_stage_inst_dmem_n4628) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2083 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5694), .Y(mem_stage_inst_dmem_n5716) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2082 ( .A(
        mem_stage_inst_dmem_ram_254__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4629) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2081 ( .A(
        mem_stage_inst_dmem_ram_254__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4630) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2080 ( .A(
        mem_stage_inst_dmem_ram_254__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4631) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2079 ( .A(
        mem_stage_inst_dmem_ram_254__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4632) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2078 ( .A(
        mem_stage_inst_dmem_ram_254__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4633) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2077 ( .A(
        mem_stage_inst_dmem_ram_254__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4634) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2076 ( .A(
        mem_stage_inst_dmem_ram_254__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4635) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2075 ( .A(
        mem_stage_inst_dmem_ram_254__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4636) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2074 ( .A(
        mem_stage_inst_dmem_ram_254__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4637) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2073 ( .A(
        mem_stage_inst_dmem_ram_254__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4638) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2072 ( .A(
        mem_stage_inst_dmem_ram_254__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4639) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2071 ( .A(
        mem_stage_inst_dmem_ram_254__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4640) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2070 ( .A(
        mem_stage_inst_dmem_ram_254__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4641) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2069 ( .A(
        mem_stage_inst_dmem_ram_254__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4642) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2068 ( .A(
        mem_stage_inst_dmem_ram_254__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4643) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2067 ( .A(
        mem_stage_inst_dmem_ram_254__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5716), .Y(mem_stage_inst_dmem_n4644) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2066 ( .A(mem_stage_inst_dmem_n5715), 
        .B(mem_stage_inst_dmem_n5691), .Y(mem_stage_inst_dmem_n5714) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2065 ( .A(
        mem_stage_inst_dmem_ram_255__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4645) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2064 ( .A(
        mem_stage_inst_dmem_ram_255__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4646) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2063 ( .A(
        mem_stage_inst_dmem_ram_255__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4647) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2062 ( .A(
        mem_stage_inst_dmem_ram_255__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4648) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2061 ( .A(
        mem_stage_inst_dmem_ram_255__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4649) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2060 ( .A(
        mem_stage_inst_dmem_ram_255__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4650) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2059 ( .A(
        mem_stage_inst_dmem_ram_255__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4651) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2058 ( .A(
        mem_stage_inst_dmem_ram_255__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4652) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2057 ( .A(
        mem_stage_inst_dmem_ram_255__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4653) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2056 ( .A(
        mem_stage_inst_dmem_ram_255__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4654) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2055 ( .A(
        mem_stage_inst_dmem_ram_255__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4655) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2054 ( .A(
        mem_stage_inst_dmem_ram_255__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4656) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2053 ( .A(
        mem_stage_inst_dmem_ram_255__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4657) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2052 ( .A(
        mem_stage_inst_dmem_ram_255__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4658) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2051 ( .A(
        mem_stage_inst_dmem_ram_255__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4659) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2050 ( .A(
        mem_stage_inst_dmem_ram_255__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5714), .Y(mem_stage_inst_dmem_n4660) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2049 ( .A(mem_stage_inst_dmem_n5712), 
        .B(mem_stage_inst_dmem_n5713), .Y(mem_stage_inst_dmem_n5692) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2048 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5689), .Y(mem_stage_inst_dmem_n5711) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2047 ( .A(
        mem_stage_inst_dmem_ram_0__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n565) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2046 ( .A(
        mem_stage_inst_dmem_ram_0__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n566) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2045 ( .A(
        mem_stage_inst_dmem_ram_0__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n567) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2044 ( .A(
        mem_stage_inst_dmem_ram_0__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n568) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2043 ( .A(
        mem_stage_inst_dmem_ram_0__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n569) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2042 ( .A(
        mem_stage_inst_dmem_ram_0__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n570) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2041 ( .A(
        mem_stage_inst_dmem_ram_0__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n571) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2040 ( .A(
        mem_stage_inst_dmem_ram_0__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n572) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2039 ( .A(
        mem_stage_inst_dmem_ram_0__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n573) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2038 ( .A(
        mem_stage_inst_dmem_ram_0__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n574) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2037 ( .A(
        mem_stage_inst_dmem_ram_0__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n575) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2036 ( .A(
        mem_stage_inst_dmem_ram_0__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n576) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2035 ( .A(
        mem_stage_inst_dmem_ram_0__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n577) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2034 ( .A(
        mem_stage_inst_dmem_ram_0__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n578) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2033 ( .A(
        mem_stage_inst_dmem_ram_0__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n579) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2032 ( .A(
        mem_stage_inst_dmem_ram_0__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5711), .Y(mem_stage_inst_dmem_n580) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2031 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5687), .Y(mem_stage_inst_dmem_n5710) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2030 ( .A(
        mem_stage_inst_dmem_ram_1__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n581) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2029 ( .A(
        mem_stage_inst_dmem_ram_1__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n582) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2028 ( .A(
        mem_stage_inst_dmem_ram_1__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n583) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2027 ( .A(
        mem_stage_inst_dmem_ram_1__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n584) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2026 ( .A(
        mem_stage_inst_dmem_ram_1__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n585) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2025 ( .A(
        mem_stage_inst_dmem_ram_1__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n586) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2024 ( .A(
        mem_stage_inst_dmem_ram_1__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n587) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2023 ( .A(
        mem_stage_inst_dmem_ram_1__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n588) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2022 ( .A(
        mem_stage_inst_dmem_ram_1__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n589) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2021 ( .A(
        mem_stage_inst_dmem_ram_1__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n590) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2020 ( .A(
        mem_stage_inst_dmem_ram_1__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n591) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2019 ( .A(
        mem_stage_inst_dmem_ram_1__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n592) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2018 ( .A(
        mem_stage_inst_dmem_ram_1__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n593) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2017 ( .A(
        mem_stage_inst_dmem_ram_1__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n594) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2016 ( .A(
        mem_stage_inst_dmem_ram_1__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n595) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2015 ( .A(
        mem_stage_inst_dmem_ram_1__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5710), .Y(mem_stage_inst_dmem_n596) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u2014 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5685), .Y(mem_stage_inst_dmem_n5709) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2013 ( .A(
        mem_stage_inst_dmem_ram_2__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n597) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2012 ( .A(
        mem_stage_inst_dmem_ram_2__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n598) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2011 ( .A(
        mem_stage_inst_dmem_ram_2__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n599) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2010 ( .A(
        mem_stage_inst_dmem_ram_2__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n600) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2009 ( .A(
        mem_stage_inst_dmem_ram_2__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n601) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2008 ( .A(
        mem_stage_inst_dmem_ram_2__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n602) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2007 ( .A(
        mem_stage_inst_dmem_ram_2__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n603) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2006 ( .A(
        mem_stage_inst_dmem_ram_2__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n604) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2005 ( .A(
        mem_stage_inst_dmem_ram_2__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n605) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2004 ( .A(
        mem_stage_inst_dmem_ram_2__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n606) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2003 ( .A(
        mem_stage_inst_dmem_ram_2__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n607) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2002 ( .A(
        mem_stage_inst_dmem_ram_2__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n608) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2001 ( .A(
        mem_stage_inst_dmem_ram_2__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n609) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u2000 ( .A(
        mem_stage_inst_dmem_ram_2__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n610) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1999 ( .A(
        mem_stage_inst_dmem_ram_2__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n611) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1998 ( .A(
        mem_stage_inst_dmem_ram_2__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5709), .Y(mem_stage_inst_dmem_n612) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1997 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5683), .Y(mem_stage_inst_dmem_n5708) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1996 ( .A(
        mem_stage_inst_dmem_ram_3__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n613) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1995 ( .A(
        mem_stage_inst_dmem_ram_3__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n614) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1994 ( .A(
        mem_stage_inst_dmem_ram_3__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n615) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1993 ( .A(
        mem_stage_inst_dmem_ram_3__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n616) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1992 ( .A(
        mem_stage_inst_dmem_ram_3__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n617) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1991 ( .A(
        mem_stage_inst_dmem_ram_3__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n618) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1990 ( .A(
        mem_stage_inst_dmem_ram_3__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n619) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1989 ( .A(
        mem_stage_inst_dmem_ram_3__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n620) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1988 ( .A(
        mem_stage_inst_dmem_ram_3__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n621) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1987 ( .A(
        mem_stage_inst_dmem_ram_3__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n622) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1986 ( .A(
        mem_stage_inst_dmem_ram_3__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n623) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1985 ( .A(
        mem_stage_inst_dmem_ram_3__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n624) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1984 ( .A(
        mem_stage_inst_dmem_ram_3__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n625) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1983 ( .A(
        mem_stage_inst_dmem_ram_3__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n626) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1982 ( .A(
        mem_stage_inst_dmem_ram_3__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n627) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1981 ( .A(
        mem_stage_inst_dmem_ram_3__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5708), .Y(mem_stage_inst_dmem_n628) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1980 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5681), .Y(mem_stage_inst_dmem_n5707) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1979 ( .A(
        mem_stage_inst_dmem_ram_4__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n629) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1978 ( .A(
        mem_stage_inst_dmem_ram_4__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n630) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1977 ( .A(
        mem_stage_inst_dmem_ram_4__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n631) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1976 ( .A(
        mem_stage_inst_dmem_ram_4__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n632) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1975 ( .A(
        mem_stage_inst_dmem_ram_4__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n633) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1974 ( .A(
        mem_stage_inst_dmem_ram_4__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n634) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1973 ( .A(
        mem_stage_inst_dmem_ram_4__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n635) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1972 ( .A(
        mem_stage_inst_dmem_ram_4__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n636) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1971 ( .A(
        mem_stage_inst_dmem_ram_4__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n637) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1970 ( .A(
        mem_stage_inst_dmem_ram_4__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n638) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1969 ( .A(
        mem_stage_inst_dmem_ram_4__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n639) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1968 ( .A(
        mem_stage_inst_dmem_ram_4__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n640) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1967 ( .A(
        mem_stage_inst_dmem_ram_4__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n641) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1966 ( .A(
        mem_stage_inst_dmem_ram_4__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n642) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1965 ( .A(
        mem_stage_inst_dmem_ram_4__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n643) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1964 ( .A(
        mem_stage_inst_dmem_ram_4__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5707), .Y(mem_stage_inst_dmem_n644) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1963 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5679), .Y(mem_stage_inst_dmem_n5706) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1962 ( .A(
        mem_stage_inst_dmem_ram_5__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n645) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1961 ( .A(
        mem_stage_inst_dmem_ram_5__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n646) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1960 ( .A(
        mem_stage_inst_dmem_ram_5__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n647) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1959 ( .A(
        mem_stage_inst_dmem_ram_5__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n648) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1958 ( .A(
        mem_stage_inst_dmem_ram_5__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n649) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1957 ( .A(
        mem_stage_inst_dmem_ram_5__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n650) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1956 ( .A(
        mem_stage_inst_dmem_ram_5__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n651) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1955 ( .A(
        mem_stage_inst_dmem_ram_5__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n652) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1954 ( .A(
        mem_stage_inst_dmem_ram_5__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n653) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1953 ( .A(
        mem_stage_inst_dmem_ram_5__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n654) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1952 ( .A(
        mem_stage_inst_dmem_ram_5__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n655) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1951 ( .A(
        mem_stage_inst_dmem_ram_5__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n656) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1950 ( .A(
        mem_stage_inst_dmem_ram_5__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n657) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1949 ( .A(
        mem_stage_inst_dmem_ram_5__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n658) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1948 ( .A(
        mem_stage_inst_dmem_ram_5__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n659) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1947 ( .A(
        mem_stage_inst_dmem_ram_5__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5706), .Y(mem_stage_inst_dmem_n660) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1946 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5677), .Y(mem_stage_inst_dmem_n5705) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1945 ( .A(
        mem_stage_inst_dmem_ram_6__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n661) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1944 ( .A(
        mem_stage_inst_dmem_ram_6__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n662) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1943 ( .A(
        mem_stage_inst_dmem_ram_6__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n663) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1942 ( .A(
        mem_stage_inst_dmem_ram_6__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n664) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1941 ( .A(
        mem_stage_inst_dmem_ram_6__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n665) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1940 ( .A(
        mem_stage_inst_dmem_ram_6__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n666) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1939 ( .A(
        mem_stage_inst_dmem_ram_6__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n667) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1938 ( .A(
        mem_stage_inst_dmem_ram_6__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n668) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1937 ( .A(
        mem_stage_inst_dmem_ram_6__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n669) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1936 ( .A(
        mem_stage_inst_dmem_ram_6__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n670) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1935 ( .A(
        mem_stage_inst_dmem_ram_6__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n671) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1934 ( .A(
        mem_stage_inst_dmem_ram_6__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n672) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1933 ( .A(
        mem_stage_inst_dmem_ram_6__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n673) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1932 ( .A(
        mem_stage_inst_dmem_ram_6__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n674) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1931 ( .A(
        mem_stage_inst_dmem_ram_6__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n675) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1930 ( .A(
        mem_stage_inst_dmem_ram_6__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5705), .Y(mem_stage_inst_dmem_n676) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1929 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5675), .Y(mem_stage_inst_dmem_n5704) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1928 ( .A(
        mem_stage_inst_dmem_ram_7__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n677) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1927 ( .A(
        mem_stage_inst_dmem_ram_7__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n678) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1926 ( .A(
        mem_stage_inst_dmem_ram_7__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n679) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1925 ( .A(
        mem_stage_inst_dmem_ram_7__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n680) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1924 ( .A(
        mem_stage_inst_dmem_ram_7__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n681) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1923 ( .A(
        mem_stage_inst_dmem_ram_7__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n682) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1922 ( .A(
        mem_stage_inst_dmem_ram_7__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n683) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1921 ( .A(
        mem_stage_inst_dmem_ram_7__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n684) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1920 ( .A(
        mem_stage_inst_dmem_ram_7__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n685) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1919 ( .A(
        mem_stage_inst_dmem_ram_7__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n686) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1918 ( .A(
        mem_stage_inst_dmem_ram_7__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n687) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1917 ( .A(
        mem_stage_inst_dmem_ram_7__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n688) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1916 ( .A(
        mem_stage_inst_dmem_ram_7__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n689) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1915 ( .A(
        mem_stage_inst_dmem_ram_7__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n690) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1914 ( .A(
        mem_stage_inst_dmem_ram_7__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n691) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1913 ( .A(
        mem_stage_inst_dmem_ram_7__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5704), .Y(mem_stage_inst_dmem_n692) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1912 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5673), .Y(mem_stage_inst_dmem_n5703) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1911 ( .A(
        mem_stage_inst_dmem_ram_8__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n693) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1910 ( .A(
        mem_stage_inst_dmem_ram_8__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n694) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1909 ( .A(
        mem_stage_inst_dmem_ram_8__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n695) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1908 ( .A(
        mem_stage_inst_dmem_ram_8__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n696) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1907 ( .A(
        mem_stage_inst_dmem_ram_8__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n697) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1906 ( .A(
        mem_stage_inst_dmem_ram_8__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n698) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1905 ( .A(
        mem_stage_inst_dmem_ram_8__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n699) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1904 ( .A(
        mem_stage_inst_dmem_ram_8__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n700) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1903 ( .A(
        mem_stage_inst_dmem_ram_8__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n701) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1902 ( .A(
        mem_stage_inst_dmem_ram_8__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n702) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1901 ( .A(
        mem_stage_inst_dmem_ram_8__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n703) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1900 ( .A(
        mem_stage_inst_dmem_ram_8__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n704) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1899 ( .A(
        mem_stage_inst_dmem_ram_8__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n705) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1898 ( .A(
        mem_stage_inst_dmem_ram_8__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n706) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1897 ( .A(
        mem_stage_inst_dmem_ram_8__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n707) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1896 ( .A(
        mem_stage_inst_dmem_ram_8__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5703), .Y(mem_stage_inst_dmem_n708) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1895 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5671), .Y(mem_stage_inst_dmem_n5702) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1894 ( .A(
        mem_stage_inst_dmem_ram_9__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n709) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1893 ( .A(
        mem_stage_inst_dmem_ram_9__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n710) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1892 ( .A(
        mem_stage_inst_dmem_ram_9__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n711) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1891 ( .A(
        mem_stage_inst_dmem_ram_9__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n712) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1890 ( .A(
        mem_stage_inst_dmem_ram_9__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n713) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1889 ( .A(
        mem_stage_inst_dmem_ram_9__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n714) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1888 ( .A(
        mem_stage_inst_dmem_ram_9__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n715) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1887 ( .A(
        mem_stage_inst_dmem_ram_9__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n716) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1886 ( .A(
        mem_stage_inst_dmem_ram_9__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n717) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1885 ( .A(
        mem_stage_inst_dmem_ram_9__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n718) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1884 ( .A(
        mem_stage_inst_dmem_ram_9__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n719) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1883 ( .A(
        mem_stage_inst_dmem_ram_9__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n720) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1882 ( .A(
        mem_stage_inst_dmem_ram_9__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n721) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1881 ( .A(
        mem_stage_inst_dmem_ram_9__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n722) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1880 ( .A(
        mem_stage_inst_dmem_ram_9__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n723) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1879 ( .A(
        mem_stage_inst_dmem_ram_9__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5702), .Y(mem_stage_inst_dmem_n724) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1878 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5668), .Y(mem_stage_inst_dmem_n5701) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1877 ( .A(
        mem_stage_inst_dmem_ram_10__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n725) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1876 ( .A(
        mem_stage_inst_dmem_ram_10__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n726) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1875 ( .A(
        mem_stage_inst_dmem_ram_10__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n727) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1874 ( .A(
        mem_stage_inst_dmem_ram_10__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n728) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1873 ( .A(
        mem_stage_inst_dmem_ram_10__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n729) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1872 ( .A(
        mem_stage_inst_dmem_ram_10__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n730) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1871 ( .A(
        mem_stage_inst_dmem_ram_10__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n731) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1870 ( .A(
        mem_stage_inst_dmem_ram_10__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n732) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1869 ( .A(
        mem_stage_inst_dmem_ram_10__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n733) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1868 ( .A(
        mem_stage_inst_dmem_ram_10__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n734) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1867 ( .A(
        mem_stage_inst_dmem_ram_10__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n735) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1866 ( .A(
        mem_stage_inst_dmem_ram_10__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n736) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1865 ( .A(
        mem_stage_inst_dmem_ram_10__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n737) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1864 ( .A(
        mem_stage_inst_dmem_ram_10__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n738) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1863 ( .A(
        mem_stage_inst_dmem_ram_10__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n739) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1862 ( .A(
        mem_stage_inst_dmem_ram_10__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5701), .Y(mem_stage_inst_dmem_n740) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1861 ( .A(mem_stage_inst_dmem_n5692), 
        .B(mem_stage_inst_dmem_n5700), .Y(mem_stage_inst_dmem_n5699) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1860 ( .A(
        mem_stage_inst_dmem_ram_11__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n741) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1859 ( .A(
        mem_stage_inst_dmem_ram_11__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n742) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1858 ( .A(
        mem_stage_inst_dmem_ram_11__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n743) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1857 ( .A(
        mem_stage_inst_dmem_ram_11__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n744) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1856 ( .A(
        mem_stage_inst_dmem_ram_11__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n745) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1855 ( .A(
        mem_stage_inst_dmem_ram_11__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n746) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1854 ( .A(
        mem_stage_inst_dmem_ram_11__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n747) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1853 ( .A(
        mem_stage_inst_dmem_ram_11__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n748) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1852 ( .A(
        mem_stage_inst_dmem_ram_11__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n749) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1851 ( .A(
        mem_stage_inst_dmem_ram_11__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n750) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1850 ( .A(
        mem_stage_inst_dmem_ram_11__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n751) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1849 ( .A(
        mem_stage_inst_dmem_ram_11__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n752) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1848 ( .A(
        mem_stage_inst_dmem_ram_11__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n753) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1847 ( .A(
        mem_stage_inst_dmem_ram_11__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n754) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1846 ( .A(
        mem_stage_inst_dmem_ram_11__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n755) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1845 ( .A(
        mem_stage_inst_dmem_ram_11__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5699), .Y(mem_stage_inst_dmem_n756) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1844 ( .A(mem_stage_inst_dmem_n5698), 
        .B(mem_stage_inst_dmem_n5692), .Y(mem_stage_inst_dmem_n5697) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1843 ( .A(
        mem_stage_inst_dmem_ram_12__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n757) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1842 ( .A(
        mem_stage_inst_dmem_ram_12__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n758) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1841 ( .A(
        mem_stage_inst_dmem_ram_12__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n759) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1840 ( .A(
        mem_stage_inst_dmem_ram_12__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n760) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1839 ( .A(
        mem_stage_inst_dmem_ram_12__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n761) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1838 ( .A(
        mem_stage_inst_dmem_ram_12__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n762) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1837 ( .A(
        mem_stage_inst_dmem_ram_12__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n763) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1836 ( .A(
        mem_stage_inst_dmem_ram_12__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n764) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1835 ( .A(
        mem_stage_inst_dmem_ram_12__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n765) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1834 ( .A(
        mem_stage_inst_dmem_ram_12__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n766) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1833 ( .A(
        mem_stage_inst_dmem_ram_12__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n767) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1832 ( .A(
        mem_stage_inst_dmem_ram_12__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n768) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1831 ( .A(
        mem_stage_inst_dmem_ram_12__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n769) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1830 ( .A(
        mem_stage_inst_dmem_ram_12__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n770) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1829 ( .A(
        mem_stage_inst_dmem_ram_12__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n771) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1828 ( .A(
        mem_stage_inst_dmem_ram_12__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5697), .Y(mem_stage_inst_dmem_n772) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1827 ( .A(mem_stage_inst_dmem_n5696), 
        .B(mem_stage_inst_dmem_n5692), .Y(mem_stage_inst_dmem_n5695) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1826 ( .A(
        mem_stage_inst_dmem_ram_13__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n773) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1825 ( .A(
        mem_stage_inst_dmem_ram_13__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n774) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1824 ( .A(
        mem_stage_inst_dmem_ram_13__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n775) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1823 ( .A(
        mem_stage_inst_dmem_ram_13__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n776) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1822 ( .A(
        mem_stage_inst_dmem_ram_13__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n777) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1821 ( .A(
        mem_stage_inst_dmem_ram_13__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n778) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1820 ( .A(
        mem_stage_inst_dmem_ram_13__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n779) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1819 ( .A(
        mem_stage_inst_dmem_ram_13__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n780) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1818 ( .A(
        mem_stage_inst_dmem_ram_13__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n781) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1817 ( .A(
        mem_stage_inst_dmem_ram_13__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n782) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1816 ( .A(
        mem_stage_inst_dmem_ram_13__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n783) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1815 ( .A(
        mem_stage_inst_dmem_ram_13__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n784) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1814 ( .A(
        mem_stage_inst_dmem_ram_13__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n785) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1813 ( .A(
        mem_stage_inst_dmem_ram_13__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n786) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1812 ( .A(
        mem_stage_inst_dmem_ram_13__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n787) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1811 ( .A(
        mem_stage_inst_dmem_ram_13__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5695), .Y(mem_stage_inst_dmem_n788) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1810 ( .A(mem_stage_inst_dmem_n5694), 
        .B(mem_stage_inst_dmem_n5692), .Y(mem_stage_inst_dmem_n5693) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1809 ( .A(
        mem_stage_inst_dmem_ram_14__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n789) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1808 ( .A(
        mem_stage_inst_dmem_ram_14__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n790) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1807 ( .A(
        mem_stage_inst_dmem_ram_14__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n791) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1806 ( .A(
        mem_stage_inst_dmem_ram_14__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n792) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1805 ( .A(
        mem_stage_inst_dmem_ram_14__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n793) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1804 ( .A(
        mem_stage_inst_dmem_ram_14__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n794) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1803 ( .A(
        mem_stage_inst_dmem_ram_14__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n795) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1802 ( .A(
        mem_stage_inst_dmem_ram_14__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n796) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1801 ( .A(
        mem_stage_inst_dmem_ram_14__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n797) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1800 ( .A(
        mem_stage_inst_dmem_ram_14__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n798) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1799 ( .A(
        mem_stage_inst_dmem_ram_14__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n799) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1798 ( .A(
        mem_stage_inst_dmem_ram_14__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n800) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1797 ( .A(
        mem_stage_inst_dmem_ram_14__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n801) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1796 ( .A(
        mem_stage_inst_dmem_ram_14__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n802) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1795 ( .A(
        mem_stage_inst_dmem_ram_14__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n803) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1794 ( .A(
        mem_stage_inst_dmem_ram_14__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5693), .Y(mem_stage_inst_dmem_n804) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1793 ( .A(mem_stage_inst_dmem_n5691), 
        .B(mem_stage_inst_dmem_n5692), .Y(mem_stage_inst_dmem_n5690) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1792 ( .A(
        mem_stage_inst_dmem_ram_15__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n805) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1791 ( .A(
        mem_stage_inst_dmem_ram_15__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n806) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1790 ( .A(
        mem_stage_inst_dmem_ram_15__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n807) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1789 ( .A(
        mem_stage_inst_dmem_ram_15__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n808) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1788 ( .A(
        mem_stage_inst_dmem_ram_15__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n809) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1787 ( .A(
        mem_stage_inst_dmem_ram_15__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n810) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1786 ( .A(
        mem_stage_inst_dmem_ram_15__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n811) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1785 ( .A(
        mem_stage_inst_dmem_ram_15__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n812) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1784 ( .A(
        mem_stage_inst_dmem_ram_15__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n813) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1783 ( .A(
        mem_stage_inst_dmem_ram_15__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n814) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1782 ( .A(
        mem_stage_inst_dmem_ram_15__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n815) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1781 ( .A(
        mem_stage_inst_dmem_ram_15__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n816) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1780 ( .A(
        mem_stage_inst_dmem_ram_15__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n817) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1779 ( .A(
        mem_stage_inst_dmem_ram_15__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n818) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1778 ( .A(
        mem_stage_inst_dmem_ram_15__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n819) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1777 ( .A(
        mem_stage_inst_dmem_ram_15__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5690), .Y(mem_stage_inst_dmem_n820) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1776 ( .A(mem_stage_inst_dmem_n5689), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5688) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1775 ( .A(
        mem_stage_inst_dmem_ram_16__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n821) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1774 ( .A(
        mem_stage_inst_dmem_ram_16__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n822) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1773 ( .A(
        mem_stage_inst_dmem_ram_16__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n823) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1772 ( .A(
        mem_stage_inst_dmem_ram_16__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n824) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1771 ( .A(
        mem_stage_inst_dmem_ram_16__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n825) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1770 ( .A(
        mem_stage_inst_dmem_ram_16__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n826) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1769 ( .A(
        mem_stage_inst_dmem_ram_16__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n827) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1768 ( .A(
        mem_stage_inst_dmem_ram_16__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n828) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1767 ( .A(
        mem_stage_inst_dmem_ram_16__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n829) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1766 ( .A(
        mem_stage_inst_dmem_ram_16__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n830) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1765 ( .A(
        mem_stage_inst_dmem_ram_16__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n831) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1764 ( .A(
        mem_stage_inst_dmem_ram_16__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n832) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1763 ( .A(
        mem_stage_inst_dmem_ram_16__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n833) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1762 ( .A(
        mem_stage_inst_dmem_ram_16__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n834) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1761 ( .A(
        mem_stage_inst_dmem_ram_16__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n835) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1760 ( .A(
        mem_stage_inst_dmem_ram_16__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5688), .Y(mem_stage_inst_dmem_n836) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1759 ( .A(mem_stage_inst_dmem_n5687), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5686) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1758 ( .A(
        mem_stage_inst_dmem_ram_17__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n837) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1757 ( .A(
        mem_stage_inst_dmem_ram_17__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n838) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1756 ( .A(
        mem_stage_inst_dmem_ram_17__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n839) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1755 ( .A(
        mem_stage_inst_dmem_ram_17__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n840) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1754 ( .A(
        mem_stage_inst_dmem_ram_17__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n841) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1753 ( .A(
        mem_stage_inst_dmem_ram_17__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n842) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1752 ( .A(
        mem_stage_inst_dmem_ram_17__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n843) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1751 ( .A(
        mem_stage_inst_dmem_ram_17__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n844) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1750 ( .A(
        mem_stage_inst_dmem_ram_17__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n845) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1749 ( .A(
        mem_stage_inst_dmem_ram_17__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n846) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1748 ( .A(
        mem_stage_inst_dmem_ram_17__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n847) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1747 ( .A(
        mem_stage_inst_dmem_ram_17__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n848) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1746 ( .A(
        mem_stage_inst_dmem_ram_17__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n849) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1745 ( .A(
        mem_stage_inst_dmem_ram_17__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n850) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1744 ( .A(
        mem_stage_inst_dmem_ram_17__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n851) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1743 ( .A(
        mem_stage_inst_dmem_ram_17__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5686), .Y(mem_stage_inst_dmem_n852) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1742 ( .A(mem_stage_inst_dmem_n5685), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5684) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1741 ( .A(
        mem_stage_inst_dmem_ram_18__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n853) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1740 ( .A(
        mem_stage_inst_dmem_ram_18__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n854) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1739 ( .A(
        mem_stage_inst_dmem_ram_18__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n855) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1738 ( .A(
        mem_stage_inst_dmem_ram_18__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n856) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1737 ( .A(
        mem_stage_inst_dmem_ram_18__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n857) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1736 ( .A(
        mem_stage_inst_dmem_ram_18__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n858) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1735 ( .A(
        mem_stage_inst_dmem_ram_18__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n859) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1734 ( .A(
        mem_stage_inst_dmem_ram_18__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n860) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1733 ( .A(
        mem_stage_inst_dmem_ram_18__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n861) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1732 ( .A(
        mem_stage_inst_dmem_ram_18__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n862) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1731 ( .A(
        mem_stage_inst_dmem_ram_18__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n863) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1730 ( .A(
        mem_stage_inst_dmem_ram_18__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n864) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1729 ( .A(
        mem_stage_inst_dmem_ram_18__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n865) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1728 ( .A(
        mem_stage_inst_dmem_ram_18__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n866) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1727 ( .A(
        mem_stage_inst_dmem_ram_18__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n867) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1726 ( .A(
        mem_stage_inst_dmem_ram_18__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5684), .Y(mem_stage_inst_dmem_n868) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1725 ( .A(mem_stage_inst_dmem_n5683), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5682) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1724 ( .A(
        mem_stage_inst_dmem_ram_19__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n869) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1723 ( .A(
        mem_stage_inst_dmem_ram_19__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n870) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1722 ( .A(
        mem_stage_inst_dmem_ram_19__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n871) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1721 ( .A(
        mem_stage_inst_dmem_ram_19__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n872) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1720 ( .A(
        mem_stage_inst_dmem_ram_19__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n873) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1719 ( .A(
        mem_stage_inst_dmem_ram_19__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n874) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1718 ( .A(
        mem_stage_inst_dmem_ram_19__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n875) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1717 ( .A(
        mem_stage_inst_dmem_ram_19__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n876) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1716 ( .A(
        mem_stage_inst_dmem_ram_19__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n877) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1715 ( .A(
        mem_stage_inst_dmem_ram_19__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n878) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1714 ( .A(
        mem_stage_inst_dmem_ram_19__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n879) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1713 ( .A(
        mem_stage_inst_dmem_ram_19__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n880) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1712 ( .A(
        mem_stage_inst_dmem_ram_19__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n881) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1711 ( .A(
        mem_stage_inst_dmem_ram_19__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n882) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1710 ( .A(
        mem_stage_inst_dmem_ram_19__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n883) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1709 ( .A(
        mem_stage_inst_dmem_ram_19__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5682), .Y(mem_stage_inst_dmem_n884) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1708 ( .A(mem_stage_inst_dmem_n5681), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5680) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1707 ( .A(
        mem_stage_inst_dmem_ram_20__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n885) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1706 ( .A(
        mem_stage_inst_dmem_ram_20__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n886) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1705 ( .A(
        mem_stage_inst_dmem_ram_20__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n887) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1704 ( .A(
        mem_stage_inst_dmem_ram_20__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n888) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1703 ( .A(
        mem_stage_inst_dmem_ram_20__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n889) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1702 ( .A(
        mem_stage_inst_dmem_ram_20__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n890) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1701 ( .A(
        mem_stage_inst_dmem_ram_20__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n891) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1700 ( .A(
        mem_stage_inst_dmem_ram_20__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n892) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1699 ( .A(
        mem_stage_inst_dmem_ram_20__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n893) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1698 ( .A(
        mem_stage_inst_dmem_ram_20__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n894) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1697 ( .A(
        mem_stage_inst_dmem_ram_20__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n895) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1696 ( .A(
        mem_stage_inst_dmem_ram_20__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n896) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1695 ( .A(
        mem_stage_inst_dmem_ram_20__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n897) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1694 ( .A(
        mem_stage_inst_dmem_ram_20__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n898) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1693 ( .A(
        mem_stage_inst_dmem_ram_20__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n899) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1692 ( .A(
        mem_stage_inst_dmem_ram_20__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5680), .Y(mem_stage_inst_dmem_n900) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1691 ( .A(mem_stage_inst_dmem_n5679), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5678) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1690 ( .A(
        mem_stage_inst_dmem_ram_21__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n901) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1689 ( .A(
        mem_stage_inst_dmem_ram_21__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n902) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1688 ( .A(
        mem_stage_inst_dmem_ram_21__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n903) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1687 ( .A(
        mem_stage_inst_dmem_ram_21__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n904) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1686 ( .A(
        mem_stage_inst_dmem_ram_21__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n905) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1685 ( .A(
        mem_stage_inst_dmem_ram_21__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n906) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1684 ( .A(
        mem_stage_inst_dmem_ram_21__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n907) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1683 ( .A(
        mem_stage_inst_dmem_ram_21__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n908) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1682 ( .A(
        mem_stage_inst_dmem_ram_21__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n909) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1681 ( .A(
        mem_stage_inst_dmem_ram_21__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n910) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1680 ( .A(
        mem_stage_inst_dmem_ram_21__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n911) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1679 ( .A(
        mem_stage_inst_dmem_ram_21__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n912) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1678 ( .A(
        mem_stage_inst_dmem_ram_21__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n913) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1677 ( .A(
        mem_stage_inst_dmem_ram_21__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n914) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1676 ( .A(
        mem_stage_inst_dmem_ram_21__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n915) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1675 ( .A(
        mem_stage_inst_dmem_ram_21__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5678), .Y(mem_stage_inst_dmem_n916) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1674 ( .A(mem_stage_inst_dmem_n5677), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5676) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1673 ( .A(
        mem_stage_inst_dmem_ram_22__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n917) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1672 ( .A(
        mem_stage_inst_dmem_ram_22__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n918) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1671 ( .A(
        mem_stage_inst_dmem_ram_22__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n919) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1670 ( .A(
        mem_stage_inst_dmem_ram_22__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n920) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1669 ( .A(
        mem_stage_inst_dmem_ram_22__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n921) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1668 ( .A(
        mem_stage_inst_dmem_ram_22__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n922) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1667 ( .A(
        mem_stage_inst_dmem_ram_22__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n923) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1666 ( .A(
        mem_stage_inst_dmem_ram_22__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n924) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1665 ( .A(
        mem_stage_inst_dmem_ram_22__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n925) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1664 ( .A(
        mem_stage_inst_dmem_ram_22__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n926) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1663 ( .A(
        mem_stage_inst_dmem_ram_22__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n927) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1662 ( .A(
        mem_stage_inst_dmem_ram_22__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n928) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1661 ( .A(
        mem_stage_inst_dmem_ram_22__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n929) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1660 ( .A(
        mem_stage_inst_dmem_ram_22__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n930) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1659 ( .A(
        mem_stage_inst_dmem_ram_22__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n931) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1658 ( .A(
        mem_stage_inst_dmem_ram_22__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5676), .Y(mem_stage_inst_dmem_n932) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1657 ( .A(mem_stage_inst_dmem_n5675), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5674) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1656 ( .A(
        mem_stage_inst_dmem_ram_23__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n933) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1655 ( .A(
        mem_stage_inst_dmem_ram_23__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n934) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1654 ( .A(
        mem_stage_inst_dmem_ram_23__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n935) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1653 ( .A(
        mem_stage_inst_dmem_ram_23__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n936) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1652 ( .A(
        mem_stage_inst_dmem_ram_23__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n937) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1651 ( .A(
        mem_stage_inst_dmem_ram_23__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n938) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1650 ( .A(
        mem_stage_inst_dmem_ram_23__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n939) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1649 ( .A(
        mem_stage_inst_dmem_ram_23__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n940) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1648 ( .A(
        mem_stage_inst_dmem_ram_23__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n941) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1647 ( .A(
        mem_stage_inst_dmem_ram_23__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n942) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1646 ( .A(
        mem_stage_inst_dmem_ram_23__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n943) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1645 ( .A(
        mem_stage_inst_dmem_ram_23__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n944) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1644 ( .A(
        mem_stage_inst_dmem_ram_23__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n945) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1643 ( .A(
        mem_stage_inst_dmem_ram_23__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n946) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1642 ( .A(
        mem_stage_inst_dmem_ram_23__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n947) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1641 ( .A(
        mem_stage_inst_dmem_ram_23__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5674), .Y(mem_stage_inst_dmem_n948) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1640 ( .A(mem_stage_inst_dmem_n5673), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5672) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1639 ( .A(
        mem_stage_inst_dmem_ram_24__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n949) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1638 ( .A(
        mem_stage_inst_dmem_ram_24__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n950) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1637 ( .A(
        mem_stage_inst_dmem_ram_24__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n951) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1636 ( .A(
        mem_stage_inst_dmem_ram_24__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n952) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1635 ( .A(
        mem_stage_inst_dmem_ram_24__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n953) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1634 ( .A(
        mem_stage_inst_dmem_ram_24__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n954) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1633 ( .A(
        mem_stage_inst_dmem_ram_24__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n955) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1632 ( .A(
        mem_stage_inst_dmem_ram_24__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n956) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1631 ( .A(
        mem_stage_inst_dmem_ram_24__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n957) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1630 ( .A(
        mem_stage_inst_dmem_ram_24__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n958) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1629 ( .A(
        mem_stage_inst_dmem_ram_24__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n959) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1628 ( .A(
        mem_stage_inst_dmem_ram_24__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n960) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1627 ( .A(
        mem_stage_inst_dmem_ram_24__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n961) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1626 ( .A(
        mem_stage_inst_dmem_ram_24__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n962) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1625 ( .A(
        mem_stage_inst_dmem_ram_24__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n963) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1624 ( .A(
        mem_stage_inst_dmem_ram_24__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5672), .Y(mem_stage_inst_dmem_n964) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1623 ( .A(mem_stage_inst_dmem_n5671), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5670) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1622 ( .A(
        mem_stage_inst_dmem_ram_25__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n965) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1621 ( .A(
        mem_stage_inst_dmem_ram_25__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n966) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1620 ( .A(
        mem_stage_inst_dmem_ram_25__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n967) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1619 ( .A(
        mem_stage_inst_dmem_ram_25__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n968) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1618 ( .A(
        mem_stage_inst_dmem_ram_25__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n969) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1617 ( .A(
        mem_stage_inst_dmem_ram_25__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n970) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1616 ( .A(
        mem_stage_inst_dmem_ram_25__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n971) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1615 ( .A(
        mem_stage_inst_dmem_ram_25__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n972) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1614 ( .A(
        mem_stage_inst_dmem_ram_25__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n973) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1613 ( .A(
        mem_stage_inst_dmem_ram_25__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n974) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1612 ( .A(
        mem_stage_inst_dmem_ram_25__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n975) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1611 ( .A(
        mem_stage_inst_dmem_ram_25__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n976) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1610 ( .A(
        mem_stage_inst_dmem_ram_25__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n977) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1609 ( .A(
        mem_stage_inst_dmem_ram_25__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n978) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1608 ( .A(
        mem_stage_inst_dmem_ram_25__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n979) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1607 ( .A(
        mem_stage_inst_dmem_ram_25__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5670), .Y(mem_stage_inst_dmem_n980) );
  AND2_X0P5M_A12TS mem_stage_inst_dmem_u1606 ( .A(mem_stage_inst_dmem_n5668), 
        .B(mem_stage_inst_dmem_n5669), .Y(mem_stage_inst_dmem_n5667) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1605 ( .A(
        mem_stage_inst_dmem_ram_26__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n981) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1604 ( .A(
        mem_stage_inst_dmem_ram_26__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n982) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1603 ( .A(
        mem_stage_inst_dmem_ram_26__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n983) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1602 ( .A(
        mem_stage_inst_dmem_ram_26__3_), .B(ex_pipeline_reg_out[8]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n984) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1601 ( .A(
        mem_stage_inst_dmem_ram_26__4_), .B(ex_pipeline_reg_out[9]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n985) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1600 ( .A(
        mem_stage_inst_dmem_ram_26__5_), .B(ex_pipeline_reg_out[10]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n986) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1599 ( .A(
        mem_stage_inst_dmem_ram_26__6_), .B(ex_pipeline_reg_out[11]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n987) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1598 ( .A(
        mem_stage_inst_dmem_ram_26__7_), .B(ex_pipeline_reg_out[12]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n988) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1597 ( .A(
        mem_stage_inst_dmem_ram_26__8_), .B(ex_pipeline_reg_out[13]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n989) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1596 ( .A(
        mem_stage_inst_dmem_ram_26__9_), .B(ex_pipeline_reg_out[14]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n990) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1595 ( .A(
        mem_stage_inst_dmem_ram_26__10_), .B(ex_pipeline_reg_out[15]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n991) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1594 ( .A(
        mem_stage_inst_dmem_ram_26__11_), .B(ex_pipeline_reg_out[16]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n992) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1593 ( .A(
        mem_stage_inst_dmem_ram_26__12_), .B(ex_pipeline_reg_out[17]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n993) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1592 ( .A(
        mem_stage_inst_dmem_ram_26__13_), .B(ex_pipeline_reg_out[18]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n994) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1591 ( .A(
        mem_stage_inst_dmem_ram_26__14_), .B(ex_pipeline_reg_out[19]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n995) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1590 ( .A(
        mem_stage_inst_dmem_ram_26__15_), .B(ex_pipeline_reg_out[20]), .S0(
        mem_stage_inst_dmem_n5667), .Y(mem_stage_inst_dmem_n996) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1589 ( .A(
        mem_stage_inst_dmem_ram_27__0_), .B(ex_pipeline_reg_out[5]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n997) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1588 ( .A(
        mem_stage_inst_dmem_ram_27__1_), .B(ex_pipeline_reg_out[6]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n998) );
  MXT2_X0P5M_A12TS mem_stage_inst_dmem_u1587 ( .A(
        mem_stage_inst_dmem_ram_27__2_), .B(ex_pipeline_reg_out[7]), .S0(
        mem_stage_inst_dmem_n5666), .Y(mem_stage_inst_dmem_n999) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1586 ( .A(
        mem_stage_inst_dmem_ram_240__15_), .B(mem_stage_inst_dmem_ram_242__15_), .C(mem_stage_inst_dmem_ram_241__15_), .D(mem_stage_inst_dmem_ram_243__15_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n59), .Y(
        mem_stage_inst_dmem_n5583) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1585 ( .A(
        mem_stage_inst_dmem_ram_244__15_), .B(mem_stage_inst_dmem_ram_246__15_), .C(mem_stage_inst_dmem_ram_245__15_), .D(mem_stage_inst_dmem_ram_247__15_), 
        .S0(mem_stage_inst_dmem_n162), .S1(mem_stage_inst_dmem_n58), .Y(
        mem_stage_inst_dmem_n5585) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1584 ( .A(
        mem_stage_inst_dmem_ram_252__15_), .B(mem_stage_inst_dmem_ram_254__15_), .C(mem_stage_inst_dmem_ram_253__15_), .D(mem_stage_inst_dmem_ram_255__15_), 
        .S0(mem_stage_inst_dmem_n161), .S1(mem_stage_inst_dmem_n63), .Y(
        mem_stage_inst_dmem_n5586) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1583 ( .A(mem_stage_inst_dmem_n5583), 
        .B(mem_stage_inst_dmem_n5584), .C(mem_stage_inst_dmem_n5585), .D(
        mem_stage_inst_dmem_n5586), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5582) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1582 ( .A(
        mem_stage_inst_dmem_ram_112__15_), .B(mem_stage_inst_dmem_ram_114__15_), .C(mem_stage_inst_dmem_ram_113__15_), .D(mem_stage_inst_dmem_ram_115__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n46), .Y(
        mem_stage_inst_dmem_n5623) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1581 ( .A(
        mem_stage_inst_dmem_ram_116__15_), .B(mem_stage_inst_dmem_ram_118__15_), .C(mem_stage_inst_dmem_ram_117__15_), .D(mem_stage_inst_dmem_ram_119__15_), 
        .S0(mem_stage_inst_dmem_n164), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n5625) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1580 ( .A(
        mem_stage_inst_dmem_ram_124__15_), .B(mem_stage_inst_dmem_ram_126__15_), .C(mem_stage_inst_dmem_ram_125__15_), .D(mem_stage_inst_dmem_ram_127__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n44), .Y(
        mem_stage_inst_dmem_n5626) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1579 ( .A(mem_stage_inst_dmem_n5623), 
        .B(mem_stage_inst_dmem_n5624), .C(mem_stage_inst_dmem_n5625), .D(
        mem_stage_inst_dmem_n5626), .S0(mem_stage_inst_dmem_n209), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5622) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1578 ( .A(
        mem_stage_inst_dmem_ram_240__14_), .B(mem_stage_inst_dmem_ram_242__14_), .C(mem_stage_inst_dmem_ram_241__14_), .D(mem_stage_inst_dmem_ram_243__14_), 
        .S0(mem_stage_inst_dmem_n115), .S1(mem_stage_inst_dmem_n47), .Y(
        mem_stage_inst_dmem_n5499) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1577 ( .A(
        mem_stage_inst_dmem_ram_244__14_), .B(mem_stage_inst_dmem_ram_246__14_), .C(mem_stage_inst_dmem_ram_245__14_), .D(mem_stage_inst_dmem_ram_247__14_), 
        .S0(mem_stage_inst_dmem_n114), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n5501) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1576 ( .A(
        mem_stage_inst_dmem_ram_252__14_), .B(mem_stage_inst_dmem_ram_254__14_), .C(mem_stage_inst_dmem_ram_253__14_), .D(mem_stage_inst_dmem_ram_255__14_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n5502) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1575 ( .A(mem_stage_inst_dmem_n5499), 
        .B(mem_stage_inst_dmem_n5500), .C(mem_stage_inst_dmem_n5501), .D(
        mem_stage_inst_dmem_n5502), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5498) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1574 ( .A(
        mem_stage_inst_dmem_ram_112__14_), .B(mem_stage_inst_dmem_ram_114__14_), .C(mem_stage_inst_dmem_ram_113__14_), .D(mem_stage_inst_dmem_ram_115__14_), 
        .S0(mem_stage_inst_dmem_n136), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5539) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1573 ( .A(
        mem_stage_inst_dmem_ram_116__14_), .B(mem_stage_inst_dmem_ram_118__14_), .C(mem_stage_inst_dmem_ram_117__14_), .D(mem_stage_inst_dmem_ram_119__14_), 
        .S0(mem_stage_inst_dmem_n132), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5541) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1572 ( .A(
        mem_stage_inst_dmem_ram_124__14_), .B(mem_stage_inst_dmem_ram_126__14_), .C(mem_stage_inst_dmem_ram_125__14_), .D(mem_stage_inst_dmem_ram_127__14_), 
        .S0(mem_stage_inst_dmem_n131), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5542) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1571 ( .A(mem_stage_inst_dmem_n5539), 
        .B(mem_stage_inst_dmem_n5540), .C(mem_stage_inst_dmem_n5541), .D(
        mem_stage_inst_dmem_n5542), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5538) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1570 ( .A(
        mem_stage_inst_dmem_ram_240__13_), .B(mem_stage_inst_dmem_ram_242__13_), .C(mem_stage_inst_dmem_ram_241__13_), .D(mem_stage_inst_dmem_ram_243__13_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n9), .Y(
        mem_stage_inst_dmem_n5415) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1569 ( .A(
        mem_stage_inst_dmem_ram_244__13_), .B(mem_stage_inst_dmem_ram_246__13_), .C(mem_stage_inst_dmem_ram_245__13_), .D(mem_stage_inst_dmem_ram_247__13_), 
        .S0(mem_stage_inst_dmem_n103), .S1(mem_stage_inst_dmem_n17), .Y(
        mem_stage_inst_dmem_n5417) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1568 ( .A(
        mem_stage_inst_dmem_ram_252__13_), .B(mem_stage_inst_dmem_ram_254__13_), .C(mem_stage_inst_dmem_ram_253__13_), .D(mem_stage_inst_dmem_ram_255__13_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n18), .Y(
        mem_stage_inst_dmem_n5418) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1567 ( .A(mem_stage_inst_dmem_n5415), 
        .B(mem_stage_inst_dmem_n5416), .C(mem_stage_inst_dmem_n5417), .D(
        mem_stage_inst_dmem_n5418), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5414) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1566 ( .A(
        mem_stage_inst_dmem_ram_112__13_), .B(mem_stage_inst_dmem_ram_114__13_), .C(mem_stage_inst_dmem_ram_113__13_), .D(mem_stage_inst_dmem_ram_115__13_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5455) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1565 ( .A(
        mem_stage_inst_dmem_ram_116__13_), .B(mem_stage_inst_dmem_ram_118__13_), .C(mem_stage_inst_dmem_ram_117__13_), .D(mem_stage_inst_dmem_ram_119__13_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5457) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1564 ( .A(
        mem_stage_inst_dmem_ram_124__13_), .B(mem_stage_inst_dmem_ram_126__13_), .C(mem_stage_inst_dmem_ram_125__13_), .D(mem_stage_inst_dmem_ram_127__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5458) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1563 ( .A(mem_stage_inst_dmem_n5455), 
        .B(mem_stage_inst_dmem_n5456), .C(mem_stage_inst_dmem_n5457), .D(
        mem_stage_inst_dmem_n5458), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5454) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1562 ( .A(
        mem_stage_inst_dmem_ram_240__12_), .B(mem_stage_inst_dmem_ram_242__12_), .C(mem_stage_inst_dmem_ram_241__12_), .D(mem_stage_inst_dmem_ram_243__12_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n54), .Y(
        mem_stage_inst_dmem_n5331) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1561 ( .A(
        mem_stage_inst_dmem_ram_244__12_), .B(mem_stage_inst_dmem_ram_246__12_), .C(mem_stage_inst_dmem_ram_245__12_), .D(mem_stage_inst_dmem_ram_247__12_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n53), .Y(
        mem_stage_inst_dmem_n5333) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1560 ( .A(
        mem_stage_inst_dmem_ram_252__12_), .B(mem_stage_inst_dmem_ram_254__12_), .C(mem_stage_inst_dmem_ram_253__12_), .D(mem_stage_inst_dmem_ram_255__12_), 
        .S0(mem_stage_inst_dmem_n102), .S1(mem_stage_inst_dmem_n10), .Y(
        mem_stage_inst_dmem_n5334) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1559 ( .A(mem_stage_inst_dmem_n5331), 
        .B(mem_stage_inst_dmem_n5332), .C(mem_stage_inst_dmem_n5333), .D(
        mem_stage_inst_dmem_n5334), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5330) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1558 ( .A(
        mem_stage_inst_dmem_ram_112__12_), .B(mem_stage_inst_dmem_ram_114__12_), .C(mem_stage_inst_dmem_ram_113__12_), .D(mem_stage_inst_dmem_ram_115__12_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5371) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1557 ( .A(
        mem_stage_inst_dmem_ram_116__12_), .B(mem_stage_inst_dmem_ram_118__12_), .C(mem_stage_inst_dmem_ram_117__12_), .D(mem_stage_inst_dmem_ram_119__12_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5373) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1556 ( .A(
        mem_stage_inst_dmem_ram_124__12_), .B(mem_stage_inst_dmem_ram_126__12_), .C(mem_stage_inst_dmem_ram_125__12_), .D(mem_stage_inst_dmem_ram_127__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5374) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1555 ( .A(mem_stage_inst_dmem_n5371), 
        .B(mem_stage_inst_dmem_n5372), .C(mem_stage_inst_dmem_n5373), .D(
        mem_stage_inst_dmem_n5374), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5370) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1554 ( .A(
        mem_stage_inst_dmem_ram_240__11_), .B(mem_stage_inst_dmem_ram_242__11_), .C(mem_stage_inst_dmem_ram_241__11_), .D(mem_stage_inst_dmem_ram_243__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5247) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1553 ( .A(
        mem_stage_inst_dmem_ram_244__11_), .B(mem_stage_inst_dmem_ram_246__11_), .C(mem_stage_inst_dmem_ram_245__11_), .D(mem_stage_inst_dmem_ram_247__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5249) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1552 ( .A(
        mem_stage_inst_dmem_ram_252__11_), .B(mem_stage_inst_dmem_ram_254__11_), .C(mem_stage_inst_dmem_ram_253__11_), .D(mem_stage_inst_dmem_ram_255__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5250) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1551 ( .A(mem_stage_inst_dmem_n5247), 
        .B(mem_stage_inst_dmem_n5248), .C(mem_stage_inst_dmem_n5249), .D(
        mem_stage_inst_dmem_n5250), .S0(mem_stage_inst_dmem_n215), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5246) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1550 ( .A(
        mem_stage_inst_dmem_ram_112__11_), .B(mem_stage_inst_dmem_ram_114__11_), .C(mem_stage_inst_dmem_ram_113__11_), .D(mem_stage_inst_dmem_ram_115__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5287) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1549 ( .A(
        mem_stage_inst_dmem_ram_116__11_), .B(mem_stage_inst_dmem_ram_118__11_), .C(mem_stage_inst_dmem_ram_117__11_), .D(mem_stage_inst_dmem_ram_119__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5289) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1548 ( .A(
        mem_stage_inst_dmem_ram_124__11_), .B(mem_stage_inst_dmem_ram_126__11_), .C(mem_stage_inst_dmem_ram_125__11_), .D(mem_stage_inst_dmem_ram_127__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5290) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1547 ( .A(mem_stage_inst_dmem_n5287), 
        .B(mem_stage_inst_dmem_n5288), .C(mem_stage_inst_dmem_n5289), .D(
        mem_stage_inst_dmem_n5290), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5286) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1546 ( .A(
        mem_stage_inst_dmem_ram_240__10_), .B(mem_stage_inst_dmem_ram_242__10_), .C(mem_stage_inst_dmem_ram_241__10_), .D(mem_stage_inst_dmem_ram_243__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5163) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1545 ( .A(
        mem_stage_inst_dmem_ram_244__10_), .B(mem_stage_inst_dmem_ram_246__10_), .C(mem_stage_inst_dmem_ram_245__10_), .D(mem_stage_inst_dmem_ram_247__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5165) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1544 ( .A(
        mem_stage_inst_dmem_ram_252__10_), .B(mem_stage_inst_dmem_ram_254__10_), .C(mem_stage_inst_dmem_ram_253__10_), .D(mem_stage_inst_dmem_ram_255__10_), 
        .S0(mem_stage_inst_dmem_n103), .S1(mem_stage_inst_dmem_n5), .Y(
        mem_stage_inst_dmem_n5166) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1543 ( .A(mem_stage_inst_dmem_n5163), 
        .B(mem_stage_inst_dmem_n5164), .C(mem_stage_inst_dmem_n5165), .D(
        mem_stage_inst_dmem_n5166), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5162) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1542 ( .A(
        mem_stage_inst_dmem_ram_112__10_), .B(mem_stage_inst_dmem_ram_114__10_), .C(mem_stage_inst_dmem_ram_113__10_), .D(mem_stage_inst_dmem_ram_115__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5203) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1541 ( .A(
        mem_stage_inst_dmem_ram_116__10_), .B(mem_stage_inst_dmem_ram_118__10_), .C(mem_stage_inst_dmem_ram_117__10_), .D(mem_stage_inst_dmem_ram_119__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5205) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1540 ( .A(
        mem_stage_inst_dmem_ram_124__10_), .B(mem_stage_inst_dmem_ram_126__10_), .C(mem_stage_inst_dmem_ram_125__10_), .D(mem_stage_inst_dmem_ram_127__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5206) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1539 ( .A(mem_stage_inst_dmem_n5203), 
        .B(mem_stage_inst_dmem_n5204), .C(mem_stage_inst_dmem_n5205), .D(
        mem_stage_inst_dmem_n5206), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5202) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1538 ( .A(
        mem_stage_inst_dmem_ram_240__9_), .B(mem_stage_inst_dmem_ram_242__9_), 
        .C(mem_stage_inst_dmem_ram_241__9_), .D(
        mem_stage_inst_dmem_ram_243__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5079) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1537 ( .A(
        mem_stage_inst_dmem_ram_244__9_), .B(mem_stage_inst_dmem_ram_246__9_), 
        .C(mem_stage_inst_dmem_ram_245__9_), .D(
        mem_stage_inst_dmem_ram_247__9_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5081) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1536 ( .A(
        mem_stage_inst_dmem_ram_252__9_), .B(mem_stage_inst_dmem_ram_254__9_), 
        .C(mem_stage_inst_dmem_ram_253__9_), .D(
        mem_stage_inst_dmem_ram_255__9_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5082) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1535 ( .A(mem_stage_inst_dmem_n5079), 
        .B(mem_stage_inst_dmem_n5080), .C(mem_stage_inst_dmem_n5081), .D(
        mem_stage_inst_dmem_n5082), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5078) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1534 ( .A(
        mem_stage_inst_dmem_ram_112__9_), .B(mem_stage_inst_dmem_ram_114__9_), 
        .C(mem_stage_inst_dmem_ram_113__9_), .D(
        mem_stage_inst_dmem_ram_115__9_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5119) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1533 ( .A(
        mem_stage_inst_dmem_ram_116__9_), .B(mem_stage_inst_dmem_ram_118__9_), 
        .C(mem_stage_inst_dmem_ram_117__9_), .D(
        mem_stage_inst_dmem_ram_119__9_), .S0(mem_stage_inst_dmem_n100), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5121) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1532 ( .A(
        mem_stage_inst_dmem_ram_124__9_), .B(mem_stage_inst_dmem_ram_126__9_), 
        .C(mem_stage_inst_dmem_ram_125__9_), .D(
        mem_stage_inst_dmem_ram_127__9_), .S0(mem_stage_inst_dmem_n99), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5122) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1531 ( .A(mem_stage_inst_dmem_n5119), 
        .B(mem_stage_inst_dmem_n5120), .C(mem_stage_inst_dmem_n5121), .D(
        mem_stage_inst_dmem_n5122), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5118) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1530 ( .A(
        mem_stage_inst_dmem_ram_240__8_), .B(mem_stage_inst_dmem_ram_242__8_), 
        .C(mem_stage_inst_dmem_ram_241__8_), .D(
        mem_stage_inst_dmem_ram_243__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n4995) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1529 ( .A(
        mem_stage_inst_dmem_ram_244__8_), .B(mem_stage_inst_dmem_ram_246__8_), 
        .C(mem_stage_inst_dmem_ram_245__8_), .D(
        mem_stage_inst_dmem_ram_247__8_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n4997) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1528 ( .A(
        mem_stage_inst_dmem_ram_252__8_), .B(mem_stage_inst_dmem_ram_254__8_), 
        .C(mem_stage_inst_dmem_ram_253__8_), .D(
        mem_stage_inst_dmem_ram_255__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4998) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1527 ( .A(mem_stage_inst_dmem_n4995), 
        .B(mem_stage_inst_dmem_n4996), .C(mem_stage_inst_dmem_n4997), .D(
        mem_stage_inst_dmem_n4998), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4994) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1526 ( .A(
        mem_stage_inst_dmem_ram_112__8_), .B(mem_stage_inst_dmem_ram_114__8_), 
        .C(mem_stage_inst_dmem_ram_113__8_), .D(
        mem_stage_inst_dmem_ram_115__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5035) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1525 ( .A(
        mem_stage_inst_dmem_ram_116__8_), .B(mem_stage_inst_dmem_ram_118__8_), 
        .C(mem_stage_inst_dmem_ram_117__8_), .D(
        mem_stage_inst_dmem_ram_119__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5037) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1524 ( .A(
        mem_stage_inst_dmem_ram_124__8_), .B(mem_stage_inst_dmem_ram_126__8_), 
        .C(mem_stage_inst_dmem_ram_125__8_), .D(
        mem_stage_inst_dmem_ram_127__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5038) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1523 ( .A(mem_stage_inst_dmem_n5035), 
        .B(mem_stage_inst_dmem_n5036), .C(mem_stage_inst_dmem_n5037), .D(
        mem_stage_inst_dmem_n5038), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5034) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1522 ( .A(
        mem_stage_inst_dmem_ram_240__7_), .B(mem_stage_inst_dmem_ram_242__7_), 
        .C(mem_stage_inst_dmem_ram_241__7_), .D(
        mem_stage_inst_dmem_ram_243__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4911) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1521 ( .A(
        mem_stage_inst_dmem_ram_244__7_), .B(mem_stage_inst_dmem_ram_246__7_), 
        .C(mem_stage_inst_dmem_ram_245__7_), .D(
        mem_stage_inst_dmem_ram_247__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4913) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1520 ( .A(
        mem_stage_inst_dmem_ram_252__7_), .B(mem_stage_inst_dmem_ram_254__7_), 
        .C(mem_stage_inst_dmem_ram_253__7_), .D(
        mem_stage_inst_dmem_ram_255__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4914) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1519 ( .A(mem_stage_inst_dmem_n4911), 
        .B(mem_stage_inst_dmem_n4912), .C(mem_stage_inst_dmem_n4913), .D(
        mem_stage_inst_dmem_n4914), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4910) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1518 ( .A(
        mem_stage_inst_dmem_ram_112__7_), .B(mem_stage_inst_dmem_ram_114__7_), 
        .C(mem_stage_inst_dmem_ram_113__7_), .D(
        mem_stage_inst_dmem_ram_115__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4951) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1517 ( .A(
        mem_stage_inst_dmem_ram_116__7_), .B(mem_stage_inst_dmem_ram_118__7_), 
        .C(mem_stage_inst_dmem_ram_117__7_), .D(
        mem_stage_inst_dmem_ram_119__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4953) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1516 ( .A(
        mem_stage_inst_dmem_ram_124__7_), .B(mem_stage_inst_dmem_ram_126__7_), 
        .C(mem_stage_inst_dmem_ram_125__7_), .D(
        mem_stage_inst_dmem_ram_127__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4954) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1515 ( .A(mem_stage_inst_dmem_n4951), 
        .B(mem_stage_inst_dmem_n4952), .C(mem_stage_inst_dmem_n4953), .D(
        mem_stage_inst_dmem_n4954), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4950) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1514 ( .A(
        mem_stage_inst_dmem_ram_240__6_), .B(mem_stage_inst_dmem_ram_242__6_), 
        .C(mem_stage_inst_dmem_ram_241__6_), .D(
        mem_stage_inst_dmem_ram_243__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4827) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1513 ( .A(
        mem_stage_inst_dmem_ram_244__6_), .B(mem_stage_inst_dmem_ram_246__6_), 
        .C(mem_stage_inst_dmem_ram_245__6_), .D(
        mem_stage_inst_dmem_ram_247__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4829) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1512 ( .A(
        mem_stage_inst_dmem_ram_252__6_), .B(mem_stage_inst_dmem_ram_254__6_), 
        .C(mem_stage_inst_dmem_ram_253__6_), .D(
        mem_stage_inst_dmem_ram_255__6_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4830) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1511 ( .A(mem_stage_inst_dmem_n4827), 
        .B(mem_stage_inst_dmem_n4828), .C(mem_stage_inst_dmem_n4829), .D(
        mem_stage_inst_dmem_n4830), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4826) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1510 ( .A(
        mem_stage_inst_dmem_ram_112__6_), .B(mem_stage_inst_dmem_ram_114__6_), 
        .C(mem_stage_inst_dmem_ram_113__6_), .D(
        mem_stage_inst_dmem_ram_115__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4867) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1509 ( .A(
        mem_stage_inst_dmem_ram_116__6_), .B(mem_stage_inst_dmem_ram_118__6_), 
        .C(mem_stage_inst_dmem_ram_117__6_), .D(
        mem_stage_inst_dmem_ram_119__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4869) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1508 ( .A(
        mem_stage_inst_dmem_ram_124__6_), .B(mem_stage_inst_dmem_ram_126__6_), 
        .C(mem_stage_inst_dmem_ram_125__6_), .D(
        mem_stage_inst_dmem_ram_127__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4870) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1507 ( .A(mem_stage_inst_dmem_n4867), 
        .B(mem_stage_inst_dmem_n4868), .C(mem_stage_inst_dmem_n4869), .D(
        mem_stage_inst_dmem_n4870), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4866) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1506 ( .A(
        mem_stage_inst_dmem_ram_240__5_), .B(mem_stage_inst_dmem_ram_242__5_), 
        .C(mem_stage_inst_dmem_ram_241__5_), .D(
        mem_stage_inst_dmem_ram_243__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4743) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1505 ( .A(
        mem_stage_inst_dmem_ram_244__5_), .B(mem_stage_inst_dmem_ram_246__5_), 
        .C(mem_stage_inst_dmem_ram_245__5_), .D(
        mem_stage_inst_dmem_ram_247__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4745) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1504 ( .A(
        mem_stage_inst_dmem_ram_252__5_), .B(mem_stage_inst_dmem_ram_254__5_), 
        .C(mem_stage_inst_dmem_ram_253__5_), .D(
        mem_stage_inst_dmem_ram_255__5_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4746) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1503 ( .A(mem_stage_inst_dmem_n4743), 
        .B(mem_stage_inst_dmem_n4744), .C(mem_stage_inst_dmem_n4745), .D(
        mem_stage_inst_dmem_n4746), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4742) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1502 ( .A(
        mem_stage_inst_dmem_ram_112__5_), .B(mem_stage_inst_dmem_ram_114__5_), 
        .C(mem_stage_inst_dmem_ram_113__5_), .D(
        mem_stage_inst_dmem_ram_115__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4783) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1501 ( .A(
        mem_stage_inst_dmem_ram_116__5_), .B(mem_stage_inst_dmem_ram_118__5_), 
        .C(mem_stage_inst_dmem_ram_117__5_), .D(
        mem_stage_inst_dmem_ram_119__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4785) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1500 ( .A(
        mem_stage_inst_dmem_ram_124__5_), .B(mem_stage_inst_dmem_ram_126__5_), 
        .C(mem_stage_inst_dmem_ram_125__5_), .D(
        mem_stage_inst_dmem_ram_127__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4786) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1499 ( .A(mem_stage_inst_dmem_n4783), 
        .B(mem_stage_inst_dmem_n4784), .C(mem_stage_inst_dmem_n4785), .D(
        mem_stage_inst_dmem_n4786), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4782) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1498 ( .A(
        mem_stage_inst_dmem_ram_240__4_), .B(mem_stage_inst_dmem_ram_242__4_), 
        .C(mem_stage_inst_dmem_ram_241__4_), .D(
        mem_stage_inst_dmem_ram_243__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n563) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1497 ( .A(
        mem_stage_inst_dmem_ram_244__4_), .B(mem_stage_inst_dmem_ram_246__4_), 
        .C(mem_stage_inst_dmem_ram_245__4_), .D(
        mem_stage_inst_dmem_ram_247__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4661) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1496 ( .A(
        mem_stage_inst_dmem_ram_252__4_), .B(mem_stage_inst_dmem_ram_254__4_), 
        .C(mem_stage_inst_dmem_ram_253__4_), .D(
        mem_stage_inst_dmem_ram_255__4_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n4662) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1495 ( .A(mem_stage_inst_dmem_n563), 
        .B(mem_stage_inst_dmem_n564), .C(mem_stage_inst_dmem_n4661), .D(
        mem_stage_inst_dmem_n4662), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n562) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1494 ( .A(
        mem_stage_inst_dmem_ram_112__4_), .B(mem_stage_inst_dmem_ram_114__4_), 
        .C(mem_stage_inst_dmem_ram_113__4_), .D(
        mem_stage_inst_dmem_ram_115__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4699) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1493 ( .A(
        mem_stage_inst_dmem_ram_116__4_), .B(mem_stage_inst_dmem_ram_118__4_), 
        .C(mem_stage_inst_dmem_ram_117__4_), .D(
        mem_stage_inst_dmem_ram_119__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4701) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1492 ( .A(
        mem_stage_inst_dmem_ram_124__4_), .B(mem_stage_inst_dmem_ram_126__4_), 
        .C(mem_stage_inst_dmem_ram_125__4_), .D(
        mem_stage_inst_dmem_ram_127__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4702) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1491 ( .A(mem_stage_inst_dmem_n4699), 
        .B(mem_stage_inst_dmem_n4700), .C(mem_stage_inst_dmem_n4701), .D(
        mem_stage_inst_dmem_n4702), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4698) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1490 ( .A(
        mem_stage_inst_dmem_ram_240__3_), .B(mem_stage_inst_dmem_ram_242__3_), 
        .C(mem_stage_inst_dmem_ram_241__3_), .D(
        mem_stage_inst_dmem_ram_243__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n479) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1489 ( .A(
        mem_stage_inst_dmem_ram_244__3_), .B(mem_stage_inst_dmem_ram_246__3_), 
        .C(mem_stage_inst_dmem_ram_245__3_), .D(
        mem_stage_inst_dmem_ram_247__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n481) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1488 ( .A(
        mem_stage_inst_dmem_ram_252__3_), .B(mem_stage_inst_dmem_ram_254__3_), 
        .C(mem_stage_inst_dmem_ram_253__3_), .D(
        mem_stage_inst_dmem_ram_255__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n482) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1487 ( .A(mem_stage_inst_dmem_n479), 
        .B(mem_stage_inst_dmem_n480), .C(mem_stage_inst_dmem_n481), .D(
        mem_stage_inst_dmem_n482), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n478) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1486 ( .A(
        mem_stage_inst_dmem_ram_112__3_), .B(mem_stage_inst_dmem_ram_114__3_), 
        .C(mem_stage_inst_dmem_ram_113__3_), .D(
        mem_stage_inst_dmem_ram_115__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n519) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1485 ( .A(
        mem_stage_inst_dmem_ram_116__3_), .B(mem_stage_inst_dmem_ram_118__3_), 
        .C(mem_stage_inst_dmem_ram_117__3_), .D(
        mem_stage_inst_dmem_ram_119__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n521) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1484 ( .A(
        mem_stage_inst_dmem_ram_124__3_), .B(mem_stage_inst_dmem_ram_126__3_), 
        .C(mem_stage_inst_dmem_ram_125__3_), .D(
        mem_stage_inst_dmem_ram_127__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n522) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1483 ( .A(mem_stage_inst_dmem_n519), 
        .B(mem_stage_inst_dmem_n520), .C(mem_stage_inst_dmem_n521), .D(
        mem_stage_inst_dmem_n522), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n518) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1482 ( .A(
        mem_stage_inst_dmem_ram_240__2_), .B(mem_stage_inst_dmem_ram_242__2_), 
        .C(mem_stage_inst_dmem_ram_241__2_), .D(
        mem_stage_inst_dmem_ram_243__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n395) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1481 ( .A(
        mem_stage_inst_dmem_ram_244__2_), .B(mem_stage_inst_dmem_ram_246__2_), 
        .C(mem_stage_inst_dmem_ram_245__2_), .D(
        mem_stage_inst_dmem_ram_247__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n397) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1480 ( .A(
        mem_stage_inst_dmem_ram_252__2_), .B(mem_stage_inst_dmem_ram_254__2_), 
        .C(mem_stage_inst_dmem_ram_253__2_), .D(
        mem_stage_inst_dmem_ram_255__2_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n398) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1479 ( .A(mem_stage_inst_dmem_n395), 
        .B(mem_stage_inst_dmem_n396), .C(mem_stage_inst_dmem_n397), .D(
        mem_stage_inst_dmem_n398), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n394) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1478 ( .A(
        mem_stage_inst_dmem_ram_112__2_), .B(mem_stage_inst_dmem_ram_114__2_), 
        .C(mem_stage_inst_dmem_ram_113__2_), .D(
        mem_stage_inst_dmem_ram_115__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n435) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1477 ( .A(
        mem_stage_inst_dmem_ram_116__2_), .B(mem_stage_inst_dmem_ram_118__2_), 
        .C(mem_stage_inst_dmem_ram_117__2_), .D(
        mem_stage_inst_dmem_ram_119__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n437) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1476 ( .A(
        mem_stage_inst_dmem_ram_124__2_), .B(mem_stage_inst_dmem_ram_126__2_), 
        .C(mem_stage_inst_dmem_ram_125__2_), .D(
        mem_stage_inst_dmem_ram_127__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n438) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1475 ( .A(mem_stage_inst_dmem_n435), 
        .B(mem_stage_inst_dmem_n436), .C(mem_stage_inst_dmem_n437), .D(
        mem_stage_inst_dmem_n438), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n434) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1474 ( .A(
        mem_stage_inst_dmem_ram_240__1_), .B(mem_stage_inst_dmem_ram_242__1_), 
        .C(mem_stage_inst_dmem_ram_241__1_), .D(
        mem_stage_inst_dmem_ram_243__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n311) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1473 ( .A(
        mem_stage_inst_dmem_ram_244__1_), .B(mem_stage_inst_dmem_ram_246__1_), 
        .C(mem_stage_inst_dmem_ram_245__1_), .D(
        mem_stage_inst_dmem_ram_247__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n313) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1472 ( .A(
        mem_stage_inst_dmem_ram_252__1_), .B(mem_stage_inst_dmem_ram_254__1_), 
        .C(mem_stage_inst_dmem_ram_253__1_), .D(
        mem_stage_inst_dmem_ram_255__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n314) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1471 ( .A(mem_stage_inst_dmem_n311), 
        .B(mem_stage_inst_dmem_n312), .C(mem_stage_inst_dmem_n313), .D(
        mem_stage_inst_dmem_n314), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n310) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1470 ( .A(
        mem_stage_inst_dmem_ram_112__1_), .B(mem_stage_inst_dmem_ram_114__1_), 
        .C(mem_stage_inst_dmem_ram_113__1_), .D(
        mem_stage_inst_dmem_ram_115__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n351) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1469 ( .A(
        mem_stage_inst_dmem_ram_116__1_), .B(mem_stage_inst_dmem_ram_118__1_), 
        .C(mem_stage_inst_dmem_ram_117__1_), .D(
        mem_stage_inst_dmem_ram_119__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n353) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1468 ( .A(
        mem_stage_inst_dmem_ram_124__1_), .B(mem_stage_inst_dmem_ram_126__1_), 
        .C(mem_stage_inst_dmem_ram_125__1_), .D(
        mem_stage_inst_dmem_ram_127__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n354) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1467 ( .A(mem_stage_inst_dmem_n351), 
        .B(mem_stage_inst_dmem_n352), .C(mem_stage_inst_dmem_n353), .D(
        mem_stage_inst_dmem_n354), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n350) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1466 ( .A(
        mem_stage_inst_dmem_ram_240__0_), .B(mem_stage_inst_dmem_ram_242__0_), 
        .C(mem_stage_inst_dmem_ram_241__0_), .D(
        mem_stage_inst_dmem_ram_243__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n227) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1465 ( .A(
        mem_stage_inst_dmem_ram_244__0_), .B(mem_stage_inst_dmem_ram_246__0_), 
        .C(mem_stage_inst_dmem_ram_245__0_), .D(
        mem_stage_inst_dmem_ram_247__0_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n229) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1464 ( .A(
        mem_stage_inst_dmem_ram_252__0_), .B(mem_stage_inst_dmem_ram_254__0_), 
        .C(mem_stage_inst_dmem_ram_253__0_), .D(
        mem_stage_inst_dmem_ram_255__0_), .S0(mem_stage_inst_dmem_n99), .S1(
        mem_stage_inst_dmem_n1), .Y(mem_stage_inst_dmem_n230) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1463 ( .A(mem_stage_inst_dmem_n227), 
        .B(mem_stage_inst_dmem_n228), .C(mem_stage_inst_dmem_n229), .D(
        mem_stage_inst_dmem_n230), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n226) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1462 ( .A(
        mem_stage_inst_dmem_ram_112__0_), .B(mem_stage_inst_dmem_ram_114__0_), 
        .C(mem_stage_inst_dmem_ram_113__0_), .D(
        mem_stage_inst_dmem_ram_115__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n267) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1461 ( .A(
        mem_stage_inst_dmem_ram_116__0_), .B(mem_stage_inst_dmem_ram_118__0_), 
        .C(mem_stage_inst_dmem_ram_117__0_), .D(
        mem_stage_inst_dmem_ram_119__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n269) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1460 ( .A(
        mem_stage_inst_dmem_ram_124__0_), .B(mem_stage_inst_dmem_ram_126__0_), 
        .C(mem_stage_inst_dmem_ram_125__0_), .D(
        mem_stage_inst_dmem_ram_127__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n270) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1459 ( .A(mem_stage_inst_dmem_n267), 
        .B(mem_stage_inst_dmem_n268), .C(mem_stage_inst_dmem_n269), .D(
        mem_stage_inst_dmem_n270), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n266) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1458 ( .A(
        mem_stage_inst_dmem_ram_60__15_), .B(mem_stage_inst_dmem_ram_62__15_), 
        .C(mem_stage_inst_dmem_ram_61__15_), .D(
        mem_stage_inst_dmem_ram_63__15_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5646) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1457 ( .A(
        mem_stage_inst_dmem_ram_28__15_), .B(mem_stage_inst_dmem_ram_30__15_), 
        .C(mem_stage_inst_dmem_ram_29__15_), .D(
        mem_stage_inst_dmem_ram_31__15_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n5656) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1456 ( .A(
        mem_stage_inst_dmem_ram_12__15_), .B(mem_stage_inst_dmem_ram_14__15_), 
        .C(mem_stage_inst_dmem_ram_13__15_), .D(
        mem_stage_inst_dmem_ram_15__15_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n5661) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1455 ( .A(
        mem_stage_inst_dmem_ram_188__15_), .B(mem_stage_inst_dmem_ram_190__15_), .C(mem_stage_inst_dmem_ram_189__15_), .D(mem_stage_inst_dmem_ram_191__15_), 
        .S0(mem_stage_inst_dmem_n120), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5606) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1454 ( .A(
        mem_stage_inst_dmem_ram_156__15_), .B(mem_stage_inst_dmem_ram_158__15_), .C(mem_stage_inst_dmem_ram_157__15_), .D(mem_stage_inst_dmem_ram_159__15_), 
        .S0(mem_stage_inst_dmem_n151), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5616) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1453 ( .A(
        mem_stage_inst_dmem_ram_140__15_), .B(mem_stage_inst_dmem_ram_142__15_), .C(mem_stage_inst_dmem_ram_141__15_), .D(mem_stage_inst_dmem_ram_143__15_), 
        .S0(mem_stage_inst_dmem_n152), .S1(mem_stage_inst_dmem_n5), .Y(
        mem_stage_inst_dmem_n5621) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1452 ( .A(
        mem_stage_inst_dmem_ram_60__14_), .B(mem_stage_inst_dmem_ram_62__14_), 
        .C(mem_stage_inst_dmem_ram_61__14_), .D(
        mem_stage_inst_dmem_ram_63__14_), .S0(mem_stage_inst_dmem_n122), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5562) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1451 ( .A(
        mem_stage_inst_dmem_ram_28__14_), .B(mem_stage_inst_dmem_ram_30__14_), 
        .C(mem_stage_inst_dmem_ram_29__14_), .D(
        mem_stage_inst_dmem_ram_31__14_), .S0(mem_stage_inst_dmem_n106), .S1(
        mem_stage_inst_dmem_n25), .Y(mem_stage_inst_dmem_n5572) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1450 ( .A(
        mem_stage_inst_dmem_ram_12__14_), .B(mem_stage_inst_dmem_ram_14__14_), 
        .C(mem_stage_inst_dmem_ram_13__14_), .D(
        mem_stage_inst_dmem_ram_15__14_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n5577) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1449 ( .A(
        mem_stage_inst_dmem_ram_188__14_), .B(mem_stage_inst_dmem_ram_190__14_), .C(mem_stage_inst_dmem_ram_189__14_), .D(mem_stage_inst_dmem_ram_191__14_), 
        .S0(mem_stage_inst_dmem_n126), .S1(mem_stage_inst_dmem_n32), .Y(
        mem_stage_inst_dmem_n5522) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1448 ( .A(
        mem_stage_inst_dmem_ram_156__14_), .B(mem_stage_inst_dmem_ram_158__14_), .C(mem_stage_inst_dmem_ram_157__14_), .D(mem_stage_inst_dmem_ram_159__14_), 
        .S0(mem_stage_inst_dmem_n109), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5532) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1447 ( .A(
        mem_stage_inst_dmem_ram_140__14_), .B(mem_stage_inst_dmem_ram_142__14_), .C(mem_stage_inst_dmem_ram_141__14_), .D(mem_stage_inst_dmem_ram_143__14_), 
        .S0(mem_stage_inst_dmem_n113), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5537) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1446 ( .A(
        mem_stage_inst_dmem_ram_60__13_), .B(mem_stage_inst_dmem_ram_62__13_), 
        .C(mem_stage_inst_dmem_ram_61__13_), .D(
        mem_stage_inst_dmem_ram_63__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5478) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1445 ( .A(
        mem_stage_inst_dmem_ram_28__13_), .B(mem_stage_inst_dmem_ram_30__13_), 
        .C(mem_stage_inst_dmem_ram_29__13_), .D(
        mem_stage_inst_dmem_ram_31__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5488) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1444 ( .A(
        mem_stage_inst_dmem_ram_12__13_), .B(mem_stage_inst_dmem_ram_14__13_), 
        .C(mem_stage_inst_dmem_ram_13__13_), .D(
        mem_stage_inst_dmem_ram_15__13_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n5493) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1443 ( .A(
        mem_stage_inst_dmem_ram_188__13_), .B(mem_stage_inst_dmem_ram_190__13_), .C(mem_stage_inst_dmem_ram_189__13_), .D(mem_stage_inst_dmem_ram_191__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n5438) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1442 ( .A(
        mem_stage_inst_dmem_ram_156__13_), .B(mem_stage_inst_dmem_ram_158__13_), .C(mem_stage_inst_dmem_ram_157__13_), .D(mem_stage_inst_dmem_ram_159__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5448) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1441 ( .A(
        mem_stage_inst_dmem_ram_140__13_), .B(mem_stage_inst_dmem_ram_142__13_), .C(mem_stage_inst_dmem_ram_141__13_), .D(mem_stage_inst_dmem_ram_143__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5453) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1440 ( .A(
        mem_stage_inst_dmem_ram_60__12_), .B(mem_stage_inst_dmem_ram_62__12_), 
        .C(mem_stage_inst_dmem_ram_61__12_), .D(
        mem_stage_inst_dmem_ram_63__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n5394) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1439 ( .A(
        mem_stage_inst_dmem_ram_28__12_), .B(mem_stage_inst_dmem_ram_30__12_), 
        .C(mem_stage_inst_dmem_ram_29__12_), .D(
        mem_stage_inst_dmem_ram_31__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n5404) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1438 ( .A(
        mem_stage_inst_dmem_ram_12__12_), .B(mem_stage_inst_dmem_ram_14__12_), 
        .C(mem_stage_inst_dmem_ram_13__12_), .D(
        mem_stage_inst_dmem_ram_15__12_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5409) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1437 ( .A(
        mem_stage_inst_dmem_ram_188__12_), .B(mem_stage_inst_dmem_ram_190__12_), .C(mem_stage_inst_dmem_ram_189__12_), .D(mem_stage_inst_dmem_ram_191__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5354) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1436 ( .A(
        mem_stage_inst_dmem_ram_156__12_), .B(mem_stage_inst_dmem_ram_158__12_), .C(mem_stage_inst_dmem_ram_157__12_), .D(mem_stage_inst_dmem_ram_159__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5364) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1435 ( .A(
        mem_stage_inst_dmem_ram_140__12_), .B(mem_stage_inst_dmem_ram_142__12_), .C(mem_stage_inst_dmem_ram_141__12_), .D(mem_stage_inst_dmem_ram_143__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5369) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1434 ( .A(
        mem_stage_inst_dmem_ram_60__11_), .B(mem_stage_inst_dmem_ram_62__11_), 
        .C(mem_stage_inst_dmem_ram_61__11_), .D(
        mem_stage_inst_dmem_ram_63__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5310) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1433 ( .A(
        mem_stage_inst_dmem_ram_28__11_), .B(mem_stage_inst_dmem_ram_30__11_), 
        .C(mem_stage_inst_dmem_ram_29__11_), .D(
        mem_stage_inst_dmem_ram_31__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5320) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1432 ( .A(
        mem_stage_inst_dmem_ram_12__11_), .B(mem_stage_inst_dmem_ram_14__11_), 
        .C(mem_stage_inst_dmem_ram_13__11_), .D(
        mem_stage_inst_dmem_ram_15__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5325) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1431 ( .A(
        mem_stage_inst_dmem_ram_188__11_), .B(mem_stage_inst_dmem_ram_190__11_), .C(mem_stage_inst_dmem_ram_189__11_), .D(mem_stage_inst_dmem_ram_191__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5270) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1430 ( .A(
        mem_stage_inst_dmem_ram_156__11_), .B(mem_stage_inst_dmem_ram_158__11_), .C(mem_stage_inst_dmem_ram_157__11_), .D(mem_stage_inst_dmem_ram_159__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5280) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1429 ( .A(
        mem_stage_inst_dmem_ram_140__11_), .B(mem_stage_inst_dmem_ram_142__11_), .C(mem_stage_inst_dmem_ram_141__11_), .D(mem_stage_inst_dmem_ram_143__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5285) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1428 ( .A(
        mem_stage_inst_dmem_ram_60__10_), .B(mem_stage_inst_dmem_ram_62__10_), 
        .C(mem_stage_inst_dmem_ram_61__10_), .D(
        mem_stage_inst_dmem_ram_63__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5226) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1427 ( .A(
        mem_stage_inst_dmem_ram_28__10_), .B(mem_stage_inst_dmem_ram_30__10_), 
        .C(mem_stage_inst_dmem_ram_29__10_), .D(
        mem_stage_inst_dmem_ram_31__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5236) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1426 ( .A(
        mem_stage_inst_dmem_ram_12__10_), .B(mem_stage_inst_dmem_ram_14__10_), 
        .C(mem_stage_inst_dmem_ram_13__10_), .D(
        mem_stage_inst_dmem_ram_15__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5241) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1425 ( .A(
        mem_stage_inst_dmem_ram_188__10_), .B(mem_stage_inst_dmem_ram_190__10_), .C(mem_stage_inst_dmem_ram_189__10_), .D(mem_stage_inst_dmem_ram_191__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5186) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1424 ( .A(
        mem_stage_inst_dmem_ram_156__10_), .B(mem_stage_inst_dmem_ram_158__10_), .C(mem_stage_inst_dmem_ram_157__10_), .D(mem_stage_inst_dmem_ram_159__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5196) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1423 ( .A(
        mem_stage_inst_dmem_ram_140__10_), .B(mem_stage_inst_dmem_ram_142__10_), .C(mem_stage_inst_dmem_ram_141__10_), .D(mem_stage_inst_dmem_ram_143__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5201) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1422 ( .A(
        mem_stage_inst_dmem_ram_60__9_), .B(mem_stage_inst_dmem_ram_62__9_), 
        .C(mem_stage_inst_dmem_ram_61__9_), .D(mem_stage_inst_dmem_ram_63__9_), 
        .S0(mem_stage_inst_dmem_n102), .S1(mem_stage_inst_dmem_n16), .Y(
        mem_stage_inst_dmem_n5142) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1421 ( .A(
        mem_stage_inst_dmem_ram_28__9_), .B(mem_stage_inst_dmem_ram_30__9_), 
        .C(mem_stage_inst_dmem_ram_29__9_), .D(mem_stage_inst_dmem_ram_31__9_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n49), .Y(
        mem_stage_inst_dmem_n5152) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1420 ( .A(
        mem_stage_inst_dmem_ram_12__9_), .B(mem_stage_inst_dmem_ram_14__9_), 
        .C(mem_stage_inst_dmem_ram_13__9_), .D(mem_stage_inst_dmem_ram_15__9_), 
        .S0(mem_stage_inst_dmem_n110), .S1(mem_stage_inst_dmem_n42), .Y(
        mem_stage_inst_dmem_n5157) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1419 ( .A(
        mem_stage_inst_dmem_ram_188__9_), .B(mem_stage_inst_dmem_ram_190__9_), 
        .C(mem_stage_inst_dmem_ram_189__9_), .D(
        mem_stage_inst_dmem_ram_191__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5102) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1418 ( .A(
        mem_stage_inst_dmem_ram_156__9_), .B(mem_stage_inst_dmem_ram_158__9_), 
        .C(mem_stage_inst_dmem_ram_157__9_), .D(
        mem_stage_inst_dmem_ram_159__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5112) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1417 ( .A(
        mem_stage_inst_dmem_ram_140__9_), .B(mem_stage_inst_dmem_ram_142__9_), 
        .C(mem_stage_inst_dmem_ram_141__9_), .D(
        mem_stage_inst_dmem_ram_143__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5117) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1416 ( .A(
        mem_stage_inst_dmem_ram_60__8_), .B(mem_stage_inst_dmem_ram_62__8_), 
        .C(mem_stage_inst_dmem_ram_61__8_), .D(mem_stage_inst_dmem_ram_63__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5058) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1415 ( .A(
        mem_stage_inst_dmem_ram_28__8_), .B(mem_stage_inst_dmem_ram_30__8_), 
        .C(mem_stage_inst_dmem_ram_29__8_), .D(mem_stage_inst_dmem_ram_31__8_), 
        .S0(mem_stage_inst_dmem_n113), .S1(mem_stage_inst_dmem_n15), .Y(
        mem_stage_inst_dmem_n5068) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1414 ( .A(
        mem_stage_inst_dmem_ram_12__8_), .B(mem_stage_inst_dmem_ram_14__8_), 
        .C(mem_stage_inst_dmem_ram_13__8_), .D(mem_stage_inst_dmem_ram_15__8_), 
        .S0(mem_stage_inst_dmem_n113), .S1(mem_stage_inst_dmem_n15), .Y(
        mem_stage_inst_dmem_n5073) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1413 ( .A(
        mem_stage_inst_dmem_ram_188__8_), .B(mem_stage_inst_dmem_ram_190__8_), 
        .C(mem_stage_inst_dmem_ram_189__8_), .D(
        mem_stage_inst_dmem_ram_191__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5018) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1412 ( .A(
        mem_stage_inst_dmem_ram_156__8_), .B(mem_stage_inst_dmem_ram_158__8_), 
        .C(mem_stage_inst_dmem_ram_157__8_), .D(
        mem_stage_inst_dmem_ram_159__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5028) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1411 ( .A(
        mem_stage_inst_dmem_ram_140__8_), .B(mem_stage_inst_dmem_ram_142__8_), 
        .C(mem_stage_inst_dmem_ram_141__8_), .D(
        mem_stage_inst_dmem_ram_143__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5033) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1410 ( .A(
        mem_stage_inst_dmem_ram_60__7_), .B(mem_stage_inst_dmem_ram_62__7_), 
        .C(mem_stage_inst_dmem_ram_61__7_), .D(mem_stage_inst_dmem_ram_63__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4974) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1409 ( .A(
        mem_stage_inst_dmem_ram_28__7_), .B(mem_stage_inst_dmem_ram_30__7_), 
        .C(mem_stage_inst_dmem_ram_29__7_), .D(mem_stage_inst_dmem_ram_31__7_), 
        .S0(mem_stage_inst_dmem_n154), .S1(mem_stage_inst_dmem_n56), .Y(
        mem_stage_inst_dmem_n4984) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1408 ( .A(
        mem_stage_inst_dmem_ram_12__7_), .B(mem_stage_inst_dmem_ram_14__7_), 
        .C(mem_stage_inst_dmem_ram_13__7_), .D(mem_stage_inst_dmem_ram_15__7_), 
        .S0(mem_stage_inst_dmem_n154), .S1(mem_stage_inst_dmem_n56), .Y(
        mem_stage_inst_dmem_n4989) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1407 ( .A(
        mem_stage_inst_dmem_ram_188__7_), .B(mem_stage_inst_dmem_ram_190__7_), 
        .C(mem_stage_inst_dmem_ram_189__7_), .D(
        mem_stage_inst_dmem_ram_191__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4934) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1406 ( .A(
        mem_stage_inst_dmem_ram_156__7_), .B(mem_stage_inst_dmem_ram_158__7_), 
        .C(mem_stage_inst_dmem_ram_157__7_), .D(
        mem_stage_inst_dmem_ram_159__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4944) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1405 ( .A(
        mem_stage_inst_dmem_ram_140__7_), .B(mem_stage_inst_dmem_ram_142__7_), 
        .C(mem_stage_inst_dmem_ram_141__7_), .D(
        mem_stage_inst_dmem_ram_143__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4949) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1404 ( .A(
        mem_stage_inst_dmem_ram_60__6_), .B(mem_stage_inst_dmem_ram_62__6_), 
        .C(mem_stage_inst_dmem_ram_61__6_), .D(mem_stage_inst_dmem_ram_63__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4890) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1403 ( .A(
        mem_stage_inst_dmem_ram_28__6_), .B(mem_stage_inst_dmem_ram_30__6_), 
        .C(mem_stage_inst_dmem_ram_29__6_), .D(mem_stage_inst_dmem_ram_31__6_), 
        .S0(mem_stage_inst_dmem_n149), .S1(mem_stage_inst_dmem_n51), .Y(
        mem_stage_inst_dmem_n4900) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1402 ( .A(
        mem_stage_inst_dmem_ram_12__6_), .B(mem_stage_inst_dmem_ram_14__6_), 
        .C(mem_stage_inst_dmem_ram_13__6_), .D(mem_stage_inst_dmem_ram_15__6_), 
        .S0(mem_stage_inst_dmem_n149), .S1(mem_stage_inst_dmem_n51), .Y(
        mem_stage_inst_dmem_n4905) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1401 ( .A(
        mem_stage_inst_dmem_ram_188__6_), .B(mem_stage_inst_dmem_ram_190__6_), 
        .C(mem_stage_inst_dmem_ram_189__6_), .D(
        mem_stage_inst_dmem_ram_191__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4850) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1400 ( .A(
        mem_stage_inst_dmem_ram_156__6_), .B(mem_stage_inst_dmem_ram_158__6_), 
        .C(mem_stage_inst_dmem_ram_157__6_), .D(
        mem_stage_inst_dmem_ram_159__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4860) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1399 ( .A(
        mem_stage_inst_dmem_ram_140__6_), .B(mem_stage_inst_dmem_ram_142__6_), 
        .C(mem_stage_inst_dmem_ram_141__6_), .D(
        mem_stage_inst_dmem_ram_143__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4865) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1398 ( .A(
        mem_stage_inst_dmem_ram_60__5_), .B(mem_stage_inst_dmem_ram_62__5_), 
        .C(mem_stage_inst_dmem_ram_61__5_), .D(mem_stage_inst_dmem_ram_63__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4806) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1397 ( .A(
        mem_stage_inst_dmem_ram_28__5_), .B(mem_stage_inst_dmem_ram_30__5_), 
        .C(mem_stage_inst_dmem_ram_29__5_), .D(mem_stage_inst_dmem_ram_31__5_), 
        .S0(mem_stage_inst_dmem_n164), .S1(ex_pipeline_reg_out[22]), .Y(
        mem_stage_inst_dmem_n4816) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1396 ( .A(
        mem_stage_inst_dmem_ram_12__5_), .B(mem_stage_inst_dmem_ram_14__5_), 
        .C(mem_stage_inst_dmem_ram_13__5_), .D(mem_stage_inst_dmem_ram_15__5_), 
        .S0(mem_stage_inst_dmem_n164), .S1(ex_pipeline_reg_out[22]), .Y(
        mem_stage_inst_dmem_n4821) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1395 ( .A(
        mem_stage_inst_dmem_ram_188__5_), .B(mem_stage_inst_dmem_ram_190__5_), 
        .C(mem_stage_inst_dmem_ram_189__5_), .D(
        mem_stage_inst_dmem_ram_191__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4766) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1394 ( .A(
        mem_stage_inst_dmem_ram_156__5_), .B(mem_stage_inst_dmem_ram_158__5_), 
        .C(mem_stage_inst_dmem_ram_157__5_), .D(
        mem_stage_inst_dmem_ram_159__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4776) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1393 ( .A(
        mem_stage_inst_dmem_ram_140__5_), .B(mem_stage_inst_dmem_ram_142__5_), 
        .C(mem_stage_inst_dmem_ram_141__5_), .D(
        mem_stage_inst_dmem_ram_143__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4781) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1392 ( .A(
        mem_stage_inst_dmem_ram_60__4_), .B(mem_stage_inst_dmem_ram_62__4_), 
        .C(mem_stage_inst_dmem_ram_61__4_), .D(mem_stage_inst_dmem_ram_63__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4722) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1391 ( .A(
        mem_stage_inst_dmem_ram_28__4_), .B(mem_stage_inst_dmem_ram_30__4_), 
        .C(mem_stage_inst_dmem_ram_29__4_), .D(mem_stage_inst_dmem_ram_31__4_), 
        .S0(mem_stage_inst_dmem_n159), .S1(mem_stage_inst_dmem_n61), .Y(
        mem_stage_inst_dmem_n4732) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1390 ( .A(
        mem_stage_inst_dmem_ram_12__4_), .B(mem_stage_inst_dmem_ram_14__4_), 
        .C(mem_stage_inst_dmem_ram_13__4_), .D(mem_stage_inst_dmem_ram_15__4_), 
        .S0(mem_stage_inst_dmem_n159), .S1(mem_stage_inst_dmem_n61), .Y(
        mem_stage_inst_dmem_n4737) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1389 ( .A(
        mem_stage_inst_dmem_ram_188__4_), .B(mem_stage_inst_dmem_ram_190__4_), 
        .C(mem_stage_inst_dmem_ram_189__4_), .D(
        mem_stage_inst_dmem_ram_191__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4682) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1388 ( .A(
        mem_stage_inst_dmem_ram_156__4_), .B(mem_stage_inst_dmem_ram_158__4_), 
        .C(mem_stage_inst_dmem_ram_157__4_), .D(
        mem_stage_inst_dmem_ram_159__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4692) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1387 ( .A(
        mem_stage_inst_dmem_ram_140__4_), .B(mem_stage_inst_dmem_ram_142__4_), 
        .C(mem_stage_inst_dmem_ram_141__4_), .D(
        mem_stage_inst_dmem_ram_143__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4697) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1386 ( .A(
        mem_stage_inst_dmem_ram_60__3_), .B(mem_stage_inst_dmem_ram_62__3_), 
        .C(mem_stage_inst_dmem_ram_61__3_), .D(mem_stage_inst_dmem_ram_63__3_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n542) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1385 ( .A(
        mem_stage_inst_dmem_ram_28__3_), .B(mem_stage_inst_dmem_ram_30__3_), 
        .C(mem_stage_inst_dmem_ram_29__3_), .D(mem_stage_inst_dmem_ram_31__3_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n552) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1384 ( .A(
        mem_stage_inst_dmem_ram_12__3_), .B(mem_stage_inst_dmem_ram_14__3_), 
        .C(mem_stage_inst_dmem_ram_13__3_), .D(mem_stage_inst_dmem_ram_15__3_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n557) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1383 ( .A(
        mem_stage_inst_dmem_ram_188__3_), .B(mem_stage_inst_dmem_ram_190__3_), 
        .C(mem_stage_inst_dmem_ram_189__3_), .D(
        mem_stage_inst_dmem_ram_191__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n502) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1382 ( .A(
        mem_stage_inst_dmem_ram_156__3_), .B(mem_stage_inst_dmem_ram_158__3_), 
        .C(mem_stage_inst_dmem_ram_157__3_), .D(
        mem_stage_inst_dmem_ram_159__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n512) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1381 ( .A(
        mem_stage_inst_dmem_ram_140__3_), .B(mem_stage_inst_dmem_ram_142__3_), 
        .C(mem_stage_inst_dmem_ram_141__3_), .D(
        mem_stage_inst_dmem_ram_143__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n517) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1380 ( .A(
        mem_stage_inst_dmem_ram_60__2_), .B(mem_stage_inst_dmem_ram_62__2_), 
        .C(mem_stage_inst_dmem_ram_61__2_), .D(mem_stage_inst_dmem_ram_63__2_), 
        .S0(mem_stage_inst_dmem_n129), .S1(mem_stage_inst_dmem_n31), .Y(
        mem_stage_inst_dmem_n458) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1379 ( .A(
        mem_stage_inst_dmem_ram_28__2_), .B(mem_stage_inst_dmem_ram_30__2_), 
        .C(mem_stage_inst_dmem_ram_29__2_), .D(mem_stage_inst_dmem_ram_31__2_), 
        .S0(mem_stage_inst_dmem_n129), .S1(mem_stage_inst_dmem_n31), .Y(
        mem_stage_inst_dmem_n468) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1378 ( .A(
        mem_stage_inst_dmem_ram_12__2_), .B(mem_stage_inst_dmem_ram_14__2_), 
        .C(mem_stage_inst_dmem_ram_13__2_), .D(mem_stage_inst_dmem_ram_15__2_), 
        .S0(mem_stage_inst_dmem_n129), .S1(mem_stage_inst_dmem_n31), .Y(
        mem_stage_inst_dmem_n473) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1377 ( .A(
        mem_stage_inst_dmem_ram_188__2_), .B(mem_stage_inst_dmem_ram_190__2_), 
        .C(mem_stage_inst_dmem_ram_189__2_), .D(
        mem_stage_inst_dmem_ram_191__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n418) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1376 ( .A(
        mem_stage_inst_dmem_ram_156__2_), .B(mem_stage_inst_dmem_ram_158__2_), 
        .C(mem_stage_inst_dmem_ram_157__2_), .D(
        mem_stage_inst_dmem_ram_159__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n428) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1375 ( .A(
        mem_stage_inst_dmem_ram_140__2_), .B(mem_stage_inst_dmem_ram_142__2_), 
        .C(mem_stage_inst_dmem_ram_141__2_), .D(
        mem_stage_inst_dmem_ram_143__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n433) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1374 ( .A(
        mem_stage_inst_dmem_ram_60__1_), .B(mem_stage_inst_dmem_ram_62__1_), 
        .C(mem_stage_inst_dmem_ram_61__1_), .D(mem_stage_inst_dmem_ram_63__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n374) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1373 ( .A(
        mem_stage_inst_dmem_ram_28__1_), .B(mem_stage_inst_dmem_ram_30__1_), 
        .C(mem_stage_inst_dmem_ram_29__1_), .D(mem_stage_inst_dmem_ram_31__1_), 
        .S0(mem_stage_inst_dmem_n144), .S1(mem_stage_inst_dmem_n46), .Y(
        mem_stage_inst_dmem_n384) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1372 ( .A(
        mem_stage_inst_dmem_ram_12__1_), .B(mem_stage_inst_dmem_ram_14__1_), 
        .C(mem_stage_inst_dmem_ram_13__1_), .D(mem_stage_inst_dmem_ram_15__1_), 
        .S0(mem_stage_inst_dmem_n144), .S1(mem_stage_inst_dmem_n46), .Y(
        mem_stage_inst_dmem_n389) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1371 ( .A(
        mem_stage_inst_dmem_ram_188__1_), .B(mem_stage_inst_dmem_ram_190__1_), 
        .C(mem_stage_inst_dmem_ram_189__1_), .D(
        mem_stage_inst_dmem_ram_191__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n334) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1370 ( .A(
        mem_stage_inst_dmem_ram_156__1_), .B(mem_stage_inst_dmem_ram_158__1_), 
        .C(mem_stage_inst_dmem_ram_157__1_), .D(
        mem_stage_inst_dmem_ram_159__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n344) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1369 ( .A(
        mem_stage_inst_dmem_ram_140__1_), .B(mem_stage_inst_dmem_ram_142__1_), 
        .C(mem_stage_inst_dmem_ram_141__1_), .D(
        mem_stage_inst_dmem_ram_143__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n349) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1368 ( .A(
        mem_stage_inst_dmem_ram_60__0_), .B(mem_stage_inst_dmem_ram_62__0_), 
        .C(mem_stage_inst_dmem_ram_61__0_), .D(mem_stage_inst_dmem_ram_63__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n290) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1367 ( .A(
        mem_stage_inst_dmem_ram_28__0_), .B(mem_stage_inst_dmem_ram_30__0_), 
        .C(mem_stage_inst_dmem_ram_29__0_), .D(mem_stage_inst_dmem_ram_31__0_), 
        .S0(mem_stage_inst_dmem_n139), .S1(mem_stage_inst_dmem_n41), .Y(
        mem_stage_inst_dmem_n300) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1366 ( .A(
        mem_stage_inst_dmem_ram_12__0_), .B(mem_stage_inst_dmem_ram_14__0_), 
        .C(mem_stage_inst_dmem_ram_13__0_), .D(mem_stage_inst_dmem_ram_15__0_), 
        .S0(mem_stage_inst_dmem_n139), .S1(mem_stage_inst_dmem_n41), .Y(
        mem_stage_inst_dmem_n305) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1365 ( .A(
        mem_stage_inst_dmem_ram_188__0_), .B(mem_stage_inst_dmem_ram_190__0_), 
        .C(mem_stage_inst_dmem_ram_189__0_), .D(
        mem_stage_inst_dmem_ram_191__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n250) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1364 ( .A(
        mem_stage_inst_dmem_ram_156__0_), .B(mem_stage_inst_dmem_ram_158__0_), 
        .C(mem_stage_inst_dmem_ram_157__0_), .D(
        mem_stage_inst_dmem_ram_159__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n260) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1363 ( .A(
        mem_stage_inst_dmem_ram_140__0_), .B(mem_stage_inst_dmem_ram_142__0_), 
        .C(mem_stage_inst_dmem_ram_141__0_), .D(
        mem_stage_inst_dmem_ram_143__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n265) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1362 ( .A(
        mem_stage_inst_dmem_ram_208__15_), .B(mem_stage_inst_dmem_ram_210__15_), .C(mem_stage_inst_dmem_ram_209__15_), .D(mem_stage_inst_dmem_ram_211__15_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n52), .Y(
        mem_stage_inst_dmem_n5593) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1361 ( .A(
        mem_stage_inst_dmem_ram_212__15_), .B(mem_stage_inst_dmem_ram_214__15_), .C(mem_stage_inst_dmem_ram_213__15_), .D(mem_stage_inst_dmem_ram_215__15_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n39), .Y(
        mem_stage_inst_dmem_n5595) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1360 ( .A(
        mem_stage_inst_dmem_ram_220__15_), .B(mem_stage_inst_dmem_ram_222__15_), .C(mem_stage_inst_dmem_ram_221__15_), .D(mem_stage_inst_dmem_ram_223__15_), 
        .S0(mem_stage_inst_dmem_n135), .S1(mem_stage_inst_dmem_n12), .Y(
        mem_stage_inst_dmem_n5596) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1359 ( .A(mem_stage_inst_dmem_n5593), 
        .B(mem_stage_inst_dmem_n5594), .C(mem_stage_inst_dmem_n5595), .D(
        mem_stage_inst_dmem_n5596), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5592) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1358 ( .A(
        mem_stage_inst_dmem_ram_80__15_), .B(mem_stage_inst_dmem_ram_82__15_), 
        .C(mem_stage_inst_dmem_ram_81__15_), .D(
        mem_stage_inst_dmem_ram_83__15_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n1), .Y(mem_stage_inst_dmem_n5633) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1357 ( .A(
        mem_stage_inst_dmem_ram_84__15_), .B(mem_stage_inst_dmem_ram_86__15_), 
        .C(mem_stage_inst_dmem_ram_85__15_), .D(
        mem_stage_inst_dmem_ram_87__15_), .S0(ex_pipeline_reg_out[23]), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5635) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1356 ( .A(
        mem_stage_inst_dmem_ram_92__15_), .B(mem_stage_inst_dmem_ram_94__15_), 
        .C(mem_stage_inst_dmem_ram_93__15_), .D(
        mem_stage_inst_dmem_ram_95__15_), .S0(ex_pipeline_reg_out[23]), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5636) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1355 ( .A(mem_stage_inst_dmem_n5633), 
        .B(mem_stage_inst_dmem_n5634), .C(mem_stage_inst_dmem_n5635), .D(
        mem_stage_inst_dmem_n5636), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5632) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1354 ( .A(
        mem_stage_inst_dmem_ram_208__14_), .B(mem_stage_inst_dmem_ram_210__14_), .C(mem_stage_inst_dmem_ram_209__14_), .D(mem_stage_inst_dmem_ram_211__14_), 
        .S0(mem_stage_inst_dmem_n129), .S1(mem_stage_inst_dmem_n38), .Y(
        mem_stage_inst_dmem_n5509) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1353 ( .A(
        mem_stage_inst_dmem_ram_212__14_), .B(mem_stage_inst_dmem_ram_214__14_), .C(mem_stage_inst_dmem_ram_213__14_), .D(mem_stage_inst_dmem_ram_215__14_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n34), .Y(
        mem_stage_inst_dmem_n5511) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1352 ( .A(
        mem_stage_inst_dmem_ram_220__14_), .B(mem_stage_inst_dmem_ram_222__14_), .C(mem_stage_inst_dmem_ram_221__14_), .D(mem_stage_inst_dmem_ram_223__14_), 
        .S0(mem_stage_inst_dmem_n127), .S1(mem_stage_inst_dmem_n33), .Y(
        mem_stage_inst_dmem_n5512) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1351 ( .A(mem_stage_inst_dmem_n5509), 
        .B(mem_stage_inst_dmem_n5510), .C(mem_stage_inst_dmem_n5511), .D(
        mem_stage_inst_dmem_n5512), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5508) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1350 ( .A(
        mem_stage_inst_dmem_ram_80__14_), .B(mem_stage_inst_dmem_ram_82__14_), 
        .C(mem_stage_inst_dmem_ram_81__14_), .D(
        mem_stage_inst_dmem_ram_83__14_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5549) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1349 ( .A(
        mem_stage_inst_dmem_ram_84__14_), .B(mem_stage_inst_dmem_ram_86__14_), 
        .C(mem_stage_inst_dmem_ram_85__14_), .D(
        mem_stage_inst_dmem_ram_87__14_), .S0(mem_stage_inst_dmem_n138), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5551) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1348 ( .A(
        mem_stage_inst_dmem_ram_92__14_), .B(mem_stage_inst_dmem_ram_94__14_), 
        .C(mem_stage_inst_dmem_ram_93__14_), .D(
        mem_stage_inst_dmem_ram_95__14_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5552) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1347 ( .A(mem_stage_inst_dmem_n5549), 
        .B(mem_stage_inst_dmem_n5550), .C(mem_stage_inst_dmem_n5551), .D(
        mem_stage_inst_dmem_n5552), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5548) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1346 ( .A(
        mem_stage_inst_dmem_ram_208__13_), .B(mem_stage_inst_dmem_ram_210__13_), .C(mem_stage_inst_dmem_ram_209__13_), .D(mem_stage_inst_dmem_ram_211__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n33), .Y(
        mem_stage_inst_dmem_n5425) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1345 ( .A(
        mem_stage_inst_dmem_ram_212__13_), .B(mem_stage_inst_dmem_ram_214__13_), .C(mem_stage_inst_dmem_ram_213__13_), .D(mem_stage_inst_dmem_ram_215__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n32), .Y(
        mem_stage_inst_dmem_n5427) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1344 ( .A(
        mem_stage_inst_dmem_ram_220__13_), .B(mem_stage_inst_dmem_ram_222__13_), .C(mem_stage_inst_dmem_ram_221__13_), .D(mem_stage_inst_dmem_ram_223__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n5428) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1343 ( .A(mem_stage_inst_dmem_n5425), 
        .B(mem_stage_inst_dmem_n5426), .C(mem_stage_inst_dmem_n5427), .D(
        mem_stage_inst_dmem_n5428), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5424) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1342 ( .A(
        mem_stage_inst_dmem_ram_80__13_), .B(mem_stage_inst_dmem_ram_82__13_), 
        .C(mem_stage_inst_dmem_ram_81__13_), .D(
        mem_stage_inst_dmem_ram_83__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n5465) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1341 ( .A(
        mem_stage_inst_dmem_ram_84__13_), .B(mem_stage_inst_dmem_ram_86__13_), 
        .C(mem_stage_inst_dmem_ram_85__13_), .D(
        mem_stage_inst_dmem_ram_87__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n5467) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1340 ( .A(
        mem_stage_inst_dmem_ram_92__13_), .B(mem_stage_inst_dmem_ram_94__13_), 
        .C(mem_stage_inst_dmem_ram_93__13_), .D(
        mem_stage_inst_dmem_ram_95__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n5468) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1339 ( .A(mem_stage_inst_dmem_n5465), 
        .B(mem_stage_inst_dmem_n5466), .C(mem_stage_inst_dmem_n5467), .D(
        mem_stage_inst_dmem_n5468), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5464) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1338 ( .A(
        mem_stage_inst_dmem_ram_208__12_), .B(mem_stage_inst_dmem_ram_210__12_), .C(mem_stage_inst_dmem_ram_209__12_), .D(mem_stage_inst_dmem_ram_211__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5341) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1337 ( .A(
        mem_stage_inst_dmem_ram_212__12_), .B(mem_stage_inst_dmem_ram_214__12_), .C(mem_stage_inst_dmem_ram_213__12_), .D(mem_stage_inst_dmem_ram_215__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5343) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1336 ( .A(
        mem_stage_inst_dmem_ram_220__12_), .B(mem_stage_inst_dmem_ram_222__12_), .C(mem_stage_inst_dmem_ram_221__12_), .D(mem_stage_inst_dmem_ram_223__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5344) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1335 ( .A(mem_stage_inst_dmem_n5341), 
        .B(mem_stage_inst_dmem_n5342), .C(mem_stage_inst_dmem_n5343), .D(
        mem_stage_inst_dmem_n5344), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5340) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1334 ( .A(
        mem_stage_inst_dmem_ram_80__12_), .B(mem_stage_inst_dmem_ram_82__12_), 
        .C(mem_stage_inst_dmem_ram_81__12_), .D(
        mem_stage_inst_dmem_ram_83__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5381) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1333 ( .A(
        mem_stage_inst_dmem_ram_84__12_), .B(mem_stage_inst_dmem_ram_86__12_), 
        .C(mem_stage_inst_dmem_ram_85__12_), .D(
        mem_stage_inst_dmem_ram_87__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5383) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1332 ( .A(
        mem_stage_inst_dmem_ram_92__12_), .B(mem_stage_inst_dmem_ram_94__12_), 
        .C(mem_stage_inst_dmem_ram_93__12_), .D(
        mem_stage_inst_dmem_ram_95__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5384) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1331 ( .A(mem_stage_inst_dmem_n5381), 
        .B(mem_stage_inst_dmem_n5382), .C(mem_stage_inst_dmem_n5383), .D(
        mem_stage_inst_dmem_n5384), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5380) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1330 ( .A(
        mem_stage_inst_dmem_ram_208__11_), .B(mem_stage_inst_dmem_ram_210__11_), .C(mem_stage_inst_dmem_ram_209__11_), .D(mem_stage_inst_dmem_ram_211__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5257) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1329 ( .A(
        mem_stage_inst_dmem_ram_212__11_), .B(mem_stage_inst_dmem_ram_214__11_), .C(mem_stage_inst_dmem_ram_213__11_), .D(mem_stage_inst_dmem_ram_215__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5259) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1328 ( .A(
        mem_stage_inst_dmem_ram_220__11_), .B(mem_stage_inst_dmem_ram_222__11_), .C(mem_stage_inst_dmem_ram_221__11_), .D(mem_stage_inst_dmem_ram_223__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5260) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1327 ( .A(mem_stage_inst_dmem_n5257), 
        .B(mem_stage_inst_dmem_n5258), .C(mem_stage_inst_dmem_n5259), .D(
        mem_stage_inst_dmem_n5260), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5256) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1326 ( .A(
        mem_stage_inst_dmem_ram_80__11_), .B(mem_stage_inst_dmem_ram_82__11_), 
        .C(mem_stage_inst_dmem_ram_81__11_), .D(
        mem_stage_inst_dmem_ram_83__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5297) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1325 ( .A(
        mem_stage_inst_dmem_ram_84__11_), .B(mem_stage_inst_dmem_ram_86__11_), 
        .C(mem_stage_inst_dmem_ram_85__11_), .D(
        mem_stage_inst_dmem_ram_87__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5299) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1324 ( .A(
        mem_stage_inst_dmem_ram_92__11_), .B(mem_stage_inst_dmem_ram_94__11_), 
        .C(mem_stage_inst_dmem_ram_93__11_), .D(
        mem_stage_inst_dmem_ram_95__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5300) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1323 ( .A(mem_stage_inst_dmem_n5297), 
        .B(mem_stage_inst_dmem_n5298), .C(mem_stage_inst_dmem_n5299), .D(
        mem_stage_inst_dmem_n5300), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5296) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1322 ( .A(
        mem_stage_inst_dmem_ram_208__10_), .B(mem_stage_inst_dmem_ram_210__10_), .C(mem_stage_inst_dmem_ram_209__10_), .D(mem_stage_inst_dmem_ram_211__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5173) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1321 ( .A(
        mem_stage_inst_dmem_ram_212__10_), .B(mem_stage_inst_dmem_ram_214__10_), .C(mem_stage_inst_dmem_ram_213__10_), .D(mem_stage_inst_dmem_ram_215__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5175) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1320 ( .A(
        mem_stage_inst_dmem_ram_220__10_), .B(mem_stage_inst_dmem_ram_222__10_), .C(mem_stage_inst_dmem_ram_221__10_), .D(mem_stage_inst_dmem_ram_223__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5176) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1319 ( .A(mem_stage_inst_dmem_n5173), 
        .B(mem_stage_inst_dmem_n5174), .C(mem_stage_inst_dmem_n5175), .D(
        mem_stage_inst_dmem_n5176), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5172) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1318 ( .A(
        mem_stage_inst_dmem_ram_80__10_), .B(mem_stage_inst_dmem_ram_82__10_), 
        .C(mem_stage_inst_dmem_ram_81__10_), .D(
        mem_stage_inst_dmem_ram_83__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5213) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1317 ( .A(
        mem_stage_inst_dmem_ram_84__10_), .B(mem_stage_inst_dmem_ram_86__10_), 
        .C(mem_stage_inst_dmem_ram_85__10_), .D(
        mem_stage_inst_dmem_ram_87__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5215) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1316 ( .A(
        mem_stage_inst_dmem_ram_92__10_), .B(mem_stage_inst_dmem_ram_94__10_), 
        .C(mem_stage_inst_dmem_ram_93__10_), .D(
        mem_stage_inst_dmem_ram_95__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5216) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1315 ( .A(mem_stage_inst_dmem_n5213), 
        .B(mem_stage_inst_dmem_n5214), .C(mem_stage_inst_dmem_n5215), .D(
        mem_stage_inst_dmem_n5216), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5212) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1314 ( .A(
        mem_stage_inst_dmem_ram_208__9_), .B(mem_stage_inst_dmem_ram_210__9_), 
        .C(mem_stage_inst_dmem_ram_209__9_), .D(
        mem_stage_inst_dmem_ram_211__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5089) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1313 ( .A(
        mem_stage_inst_dmem_ram_212__9_), .B(mem_stage_inst_dmem_ram_214__9_), 
        .C(mem_stage_inst_dmem_ram_213__9_), .D(
        mem_stage_inst_dmem_ram_215__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5091) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1312 ( .A(
        mem_stage_inst_dmem_ram_220__9_), .B(mem_stage_inst_dmem_ram_222__9_), 
        .C(mem_stage_inst_dmem_ram_221__9_), .D(
        mem_stage_inst_dmem_ram_223__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5092) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1311 ( .A(mem_stage_inst_dmem_n5089), 
        .B(mem_stage_inst_dmem_n5090), .C(mem_stage_inst_dmem_n5091), .D(
        mem_stage_inst_dmem_n5092), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5088) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1310 ( .A(
        mem_stage_inst_dmem_ram_80__9_), .B(mem_stage_inst_dmem_ram_82__9_), 
        .C(mem_stage_inst_dmem_ram_81__9_), .D(mem_stage_inst_dmem_ram_83__9_), 
        .S0(mem_stage_inst_dmem_n141), .S1(mem_stage_inst_dmem_n29), .Y(
        mem_stage_inst_dmem_n5129) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1309 ( .A(
        mem_stage_inst_dmem_ram_84__9_), .B(mem_stage_inst_dmem_ram_86__9_), 
        .C(mem_stage_inst_dmem_ram_85__9_), .D(mem_stage_inst_dmem_ram_87__9_), 
        .S0(mem_stage_inst_dmem_n140), .S1(mem_stage_inst_dmem_n28), .Y(
        mem_stage_inst_dmem_n5131) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1308 ( .A(
        mem_stage_inst_dmem_ram_92__9_), .B(mem_stage_inst_dmem_ram_94__9_), 
        .C(mem_stage_inst_dmem_ram_93__9_), .D(mem_stage_inst_dmem_ram_95__9_), 
        .S0(mem_stage_inst_dmem_n159), .S1(mem_stage_inst_dmem_n18), .Y(
        mem_stage_inst_dmem_n5132) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1307 ( .A(mem_stage_inst_dmem_n5129), 
        .B(mem_stage_inst_dmem_n5130), .C(mem_stage_inst_dmem_n5131), .D(
        mem_stage_inst_dmem_n5132), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5128) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1306 ( .A(
        mem_stage_inst_dmem_ram_208__8_), .B(mem_stage_inst_dmem_ram_210__8_), 
        .C(mem_stage_inst_dmem_ram_209__8_), .D(
        mem_stage_inst_dmem_ram_211__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5005) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1305 ( .A(
        mem_stage_inst_dmem_ram_212__8_), .B(mem_stage_inst_dmem_ram_214__8_), 
        .C(mem_stage_inst_dmem_ram_213__8_), .D(
        mem_stage_inst_dmem_ram_215__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5007) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1304 ( .A(
        mem_stage_inst_dmem_ram_220__8_), .B(mem_stage_inst_dmem_ram_222__8_), 
        .C(mem_stage_inst_dmem_ram_221__8_), .D(
        mem_stage_inst_dmem_ram_223__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5008) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1303 ( .A(mem_stage_inst_dmem_n5005), 
        .B(mem_stage_inst_dmem_n5006), .C(mem_stage_inst_dmem_n5007), .D(
        mem_stage_inst_dmem_n5008), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5004) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1302 ( .A(
        mem_stage_inst_dmem_ram_80__8_), .B(mem_stage_inst_dmem_ram_82__8_), 
        .C(mem_stage_inst_dmem_ram_81__8_), .D(mem_stage_inst_dmem_ram_83__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5045) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1301 ( .A(
        mem_stage_inst_dmem_ram_84__8_), .B(mem_stage_inst_dmem_ram_86__8_), 
        .C(mem_stage_inst_dmem_ram_85__8_), .D(mem_stage_inst_dmem_ram_87__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5047) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1300 ( .A(
        mem_stage_inst_dmem_ram_92__8_), .B(mem_stage_inst_dmem_ram_94__8_), 
        .C(mem_stage_inst_dmem_ram_93__8_), .D(mem_stage_inst_dmem_ram_95__8_), 
        .S0(mem_stage_inst_dmem_n111), .S1(mem_stage_inst_dmem_n13), .Y(
        mem_stage_inst_dmem_n5048) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1299 ( .A(mem_stage_inst_dmem_n5045), 
        .B(mem_stage_inst_dmem_n5046), .C(mem_stage_inst_dmem_n5047), .D(
        mem_stage_inst_dmem_n5048), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5044) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1298 ( .A(
        mem_stage_inst_dmem_ram_208__7_), .B(mem_stage_inst_dmem_ram_210__7_), 
        .C(mem_stage_inst_dmem_ram_209__7_), .D(
        mem_stage_inst_dmem_ram_211__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4921) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1297 ( .A(
        mem_stage_inst_dmem_ram_212__7_), .B(mem_stage_inst_dmem_ram_214__7_), 
        .C(mem_stage_inst_dmem_ram_213__7_), .D(
        mem_stage_inst_dmem_ram_215__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4923) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1296 ( .A(
        mem_stage_inst_dmem_ram_220__7_), .B(mem_stage_inst_dmem_ram_222__7_), 
        .C(mem_stage_inst_dmem_ram_221__7_), .D(
        mem_stage_inst_dmem_ram_223__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4924) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1295 ( .A(mem_stage_inst_dmem_n4921), 
        .B(mem_stage_inst_dmem_n4922), .C(mem_stage_inst_dmem_n4923), .D(
        mem_stage_inst_dmem_n4924), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4920) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1294 ( .A(
        mem_stage_inst_dmem_ram_80__7_), .B(mem_stage_inst_dmem_ram_82__7_), 
        .C(mem_stage_inst_dmem_ram_81__7_), .D(mem_stage_inst_dmem_ram_83__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4961) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1293 ( .A(
        mem_stage_inst_dmem_ram_84__7_), .B(mem_stage_inst_dmem_ram_86__7_), 
        .C(mem_stage_inst_dmem_ram_85__7_), .D(mem_stage_inst_dmem_ram_87__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4963) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1292 ( .A(
        mem_stage_inst_dmem_ram_92__7_), .B(mem_stage_inst_dmem_ram_94__7_), 
        .C(mem_stage_inst_dmem_ram_93__7_), .D(mem_stage_inst_dmem_ram_95__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4964) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1291 ( .A(mem_stage_inst_dmem_n4961), 
        .B(mem_stage_inst_dmem_n4962), .C(mem_stage_inst_dmem_n4963), .D(
        mem_stage_inst_dmem_n4964), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4960) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1290 ( .A(
        mem_stage_inst_dmem_ram_208__6_), .B(mem_stage_inst_dmem_ram_210__6_), 
        .C(mem_stage_inst_dmem_ram_209__6_), .D(
        mem_stage_inst_dmem_ram_211__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4837) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1289 ( .A(
        mem_stage_inst_dmem_ram_212__6_), .B(mem_stage_inst_dmem_ram_214__6_), 
        .C(mem_stage_inst_dmem_ram_213__6_), .D(
        mem_stage_inst_dmem_ram_215__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4839) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1288 ( .A(
        mem_stage_inst_dmem_ram_220__6_), .B(mem_stage_inst_dmem_ram_222__6_), 
        .C(mem_stage_inst_dmem_ram_221__6_), .D(
        mem_stage_inst_dmem_ram_223__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4840) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1287 ( .A(mem_stage_inst_dmem_n4837), 
        .B(mem_stage_inst_dmem_n4838), .C(mem_stage_inst_dmem_n4839), .D(
        mem_stage_inst_dmem_n4840), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4836) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1286 ( .A(
        mem_stage_inst_dmem_ram_80__6_), .B(mem_stage_inst_dmem_ram_82__6_), 
        .C(mem_stage_inst_dmem_ram_81__6_), .D(mem_stage_inst_dmem_ram_83__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4877) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1285 ( .A(
        mem_stage_inst_dmem_ram_84__6_), .B(mem_stage_inst_dmem_ram_86__6_), 
        .C(mem_stage_inst_dmem_ram_85__6_), .D(mem_stage_inst_dmem_ram_87__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4879) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1284 ( .A(
        mem_stage_inst_dmem_ram_92__6_), .B(mem_stage_inst_dmem_ram_94__6_), 
        .C(mem_stage_inst_dmem_ram_93__6_), .D(mem_stage_inst_dmem_ram_95__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4880) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1283 ( .A(mem_stage_inst_dmem_n4877), 
        .B(mem_stage_inst_dmem_n4878), .C(mem_stage_inst_dmem_n4879), .D(
        mem_stage_inst_dmem_n4880), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4876) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1282 ( .A(
        mem_stage_inst_dmem_ram_208__5_), .B(mem_stage_inst_dmem_ram_210__5_), 
        .C(mem_stage_inst_dmem_ram_209__5_), .D(
        mem_stage_inst_dmem_ram_211__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4753) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1281 ( .A(
        mem_stage_inst_dmem_ram_212__5_), .B(mem_stage_inst_dmem_ram_214__5_), 
        .C(mem_stage_inst_dmem_ram_213__5_), .D(
        mem_stage_inst_dmem_ram_215__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4755) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1280 ( .A(
        mem_stage_inst_dmem_ram_220__5_), .B(mem_stage_inst_dmem_ram_222__5_), 
        .C(mem_stage_inst_dmem_ram_221__5_), .D(
        mem_stage_inst_dmem_ram_223__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4756) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1279 ( .A(mem_stage_inst_dmem_n4753), 
        .B(mem_stage_inst_dmem_n4754), .C(mem_stage_inst_dmem_n4755), .D(
        mem_stage_inst_dmem_n4756), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4752) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1278 ( .A(
        mem_stage_inst_dmem_ram_80__5_), .B(mem_stage_inst_dmem_ram_82__5_), 
        .C(mem_stage_inst_dmem_ram_81__5_), .D(mem_stage_inst_dmem_ram_83__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4793) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1277 ( .A(
        mem_stage_inst_dmem_ram_84__5_), .B(mem_stage_inst_dmem_ram_86__5_), 
        .C(mem_stage_inst_dmem_ram_85__5_), .D(mem_stage_inst_dmem_ram_87__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4795) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1276 ( .A(
        mem_stage_inst_dmem_ram_92__5_), .B(mem_stage_inst_dmem_ram_94__5_), 
        .C(mem_stage_inst_dmem_ram_93__5_), .D(mem_stage_inst_dmem_ram_95__5_), 
        .S0(mem_stage_inst_dmem_n162), .S1(mem_stage_inst_dmem_n64), .Y(
        mem_stage_inst_dmem_n4796) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1275 ( .A(mem_stage_inst_dmem_n4793), 
        .B(mem_stage_inst_dmem_n4794), .C(mem_stage_inst_dmem_n4795), .D(
        mem_stage_inst_dmem_n4796), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4792) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1274 ( .A(
        mem_stage_inst_dmem_ram_208__4_), .B(mem_stage_inst_dmem_ram_210__4_), 
        .C(mem_stage_inst_dmem_ram_209__4_), .D(
        mem_stage_inst_dmem_ram_211__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4669) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1273 ( .A(
        mem_stage_inst_dmem_ram_212__4_), .B(mem_stage_inst_dmem_ram_214__4_), 
        .C(mem_stage_inst_dmem_ram_213__4_), .D(
        mem_stage_inst_dmem_ram_215__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4671) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1272 ( .A(
        mem_stage_inst_dmem_ram_220__4_), .B(mem_stage_inst_dmem_ram_222__4_), 
        .C(mem_stage_inst_dmem_ram_221__4_), .D(
        mem_stage_inst_dmem_ram_223__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4672) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1271 ( .A(mem_stage_inst_dmem_n4669), 
        .B(mem_stage_inst_dmem_n4670), .C(mem_stage_inst_dmem_n4671), .D(
        mem_stage_inst_dmem_n4672), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4668) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1270 ( .A(
        mem_stage_inst_dmem_ram_80__4_), .B(mem_stage_inst_dmem_ram_82__4_), 
        .C(mem_stage_inst_dmem_ram_81__4_), .D(mem_stage_inst_dmem_ram_83__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4709) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1269 ( .A(
        mem_stage_inst_dmem_ram_84__4_), .B(mem_stage_inst_dmem_ram_86__4_), 
        .C(mem_stage_inst_dmem_ram_85__4_), .D(mem_stage_inst_dmem_ram_87__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4711) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1268 ( .A(
        mem_stage_inst_dmem_ram_92__4_), .B(mem_stage_inst_dmem_ram_94__4_), 
        .C(mem_stage_inst_dmem_ram_93__4_), .D(mem_stage_inst_dmem_ram_95__4_), 
        .S0(mem_stage_inst_dmem_n157), .S1(mem_stage_inst_dmem_n59), .Y(
        mem_stage_inst_dmem_n4712) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1267 ( .A(mem_stage_inst_dmem_n4709), 
        .B(mem_stage_inst_dmem_n4710), .C(mem_stage_inst_dmem_n4711), .D(
        mem_stage_inst_dmem_n4712), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4708) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1266 ( .A(
        mem_stage_inst_dmem_ram_208__3_), .B(mem_stage_inst_dmem_ram_210__3_), 
        .C(mem_stage_inst_dmem_ram_209__3_), .D(
        mem_stage_inst_dmem_ram_211__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n489) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1265 ( .A(
        mem_stage_inst_dmem_ram_212__3_), .B(mem_stage_inst_dmem_ram_214__3_), 
        .C(mem_stage_inst_dmem_ram_213__3_), .D(
        mem_stage_inst_dmem_ram_215__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n491) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1264 ( .A(
        mem_stage_inst_dmem_ram_220__3_), .B(mem_stage_inst_dmem_ram_222__3_), 
        .C(mem_stage_inst_dmem_ram_221__3_), .D(
        mem_stage_inst_dmem_ram_223__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n492) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1263 ( .A(mem_stage_inst_dmem_n489), 
        .B(mem_stage_inst_dmem_n490), .C(mem_stage_inst_dmem_n491), .D(
        mem_stage_inst_dmem_n492), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n488) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1262 ( .A(
        mem_stage_inst_dmem_ram_80__3_), .B(mem_stage_inst_dmem_ram_82__3_), 
        .C(mem_stage_inst_dmem_ram_81__3_), .D(mem_stage_inst_dmem_ram_83__3_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n529) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1261 ( .A(
        mem_stage_inst_dmem_ram_84__3_), .B(mem_stage_inst_dmem_ram_86__3_), 
        .C(mem_stage_inst_dmem_ram_85__3_), .D(mem_stage_inst_dmem_ram_87__3_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n531) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1260 ( .A(
        mem_stage_inst_dmem_ram_92__3_), .B(mem_stage_inst_dmem_ram_94__3_), 
        .C(mem_stage_inst_dmem_ram_93__3_), .D(mem_stage_inst_dmem_ram_95__3_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n532) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1259 ( .A(mem_stage_inst_dmem_n529), 
        .B(mem_stage_inst_dmem_n530), .C(mem_stage_inst_dmem_n531), .D(
        mem_stage_inst_dmem_n532), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n528) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1258 ( .A(
        mem_stage_inst_dmem_ram_208__2_), .B(mem_stage_inst_dmem_ram_210__2_), 
        .C(mem_stage_inst_dmem_ram_209__2_), .D(
        mem_stage_inst_dmem_ram_211__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n405) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1257 ( .A(
        mem_stage_inst_dmem_ram_212__2_), .B(mem_stage_inst_dmem_ram_214__2_), 
        .C(mem_stage_inst_dmem_ram_213__2_), .D(
        mem_stage_inst_dmem_ram_215__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n407) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1256 ( .A(
        mem_stage_inst_dmem_ram_220__2_), .B(mem_stage_inst_dmem_ram_222__2_), 
        .C(mem_stage_inst_dmem_ram_221__2_), .D(
        mem_stage_inst_dmem_ram_223__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n408) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1255 ( .A(mem_stage_inst_dmem_n405), 
        .B(mem_stage_inst_dmem_n406), .C(mem_stage_inst_dmem_n407), .D(
        mem_stage_inst_dmem_n408), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n404) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1254 ( .A(
        mem_stage_inst_dmem_ram_80__2_), .B(mem_stage_inst_dmem_ram_82__2_), 
        .C(mem_stage_inst_dmem_ram_81__2_), .D(mem_stage_inst_dmem_ram_83__2_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n445) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1253 ( .A(
        mem_stage_inst_dmem_ram_84__2_), .B(mem_stage_inst_dmem_ram_86__2_), 
        .C(mem_stage_inst_dmem_ram_85__2_), .D(mem_stage_inst_dmem_ram_87__2_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n447) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1252 ( .A(
        mem_stage_inst_dmem_ram_92__2_), .B(mem_stage_inst_dmem_ram_94__2_), 
        .C(mem_stage_inst_dmem_ram_93__2_), .D(mem_stage_inst_dmem_ram_95__2_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n448) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1251 ( .A(mem_stage_inst_dmem_n445), 
        .B(mem_stage_inst_dmem_n446), .C(mem_stage_inst_dmem_n447), .D(
        mem_stage_inst_dmem_n448), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n444) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1250 ( .A(
        mem_stage_inst_dmem_ram_208__1_), .B(mem_stage_inst_dmem_ram_210__1_), 
        .C(mem_stage_inst_dmem_ram_209__1_), .D(
        mem_stage_inst_dmem_ram_211__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n321) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1249 ( .A(
        mem_stage_inst_dmem_ram_212__1_), .B(mem_stage_inst_dmem_ram_214__1_), 
        .C(mem_stage_inst_dmem_ram_213__1_), .D(
        mem_stage_inst_dmem_ram_215__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n323) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1248 ( .A(
        mem_stage_inst_dmem_ram_220__1_), .B(mem_stage_inst_dmem_ram_222__1_), 
        .C(mem_stage_inst_dmem_ram_221__1_), .D(
        mem_stage_inst_dmem_ram_223__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n324) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1247 ( .A(mem_stage_inst_dmem_n321), 
        .B(mem_stage_inst_dmem_n322), .C(mem_stage_inst_dmem_n323), .D(
        mem_stage_inst_dmem_n324), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n320) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1246 ( .A(
        mem_stage_inst_dmem_ram_80__1_), .B(mem_stage_inst_dmem_ram_82__1_), 
        .C(mem_stage_inst_dmem_ram_81__1_), .D(mem_stage_inst_dmem_ram_83__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n361) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1245 ( .A(
        mem_stage_inst_dmem_ram_84__1_), .B(mem_stage_inst_dmem_ram_86__1_), 
        .C(mem_stage_inst_dmem_ram_85__1_), .D(mem_stage_inst_dmem_ram_87__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n363) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1244 ( .A(
        mem_stage_inst_dmem_ram_92__1_), .B(mem_stage_inst_dmem_ram_94__1_), 
        .C(mem_stage_inst_dmem_ram_93__1_), .D(mem_stage_inst_dmem_ram_95__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n364) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1243 ( .A(mem_stage_inst_dmem_n361), 
        .B(mem_stage_inst_dmem_n362), .C(mem_stage_inst_dmem_n363), .D(
        mem_stage_inst_dmem_n364), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n360) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1242 ( .A(
        mem_stage_inst_dmem_ram_208__0_), .B(mem_stage_inst_dmem_ram_210__0_), 
        .C(mem_stage_inst_dmem_ram_209__0_), .D(
        mem_stage_inst_dmem_ram_211__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n237) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1241 ( .A(
        mem_stage_inst_dmem_ram_212__0_), .B(mem_stage_inst_dmem_ram_214__0_), 
        .C(mem_stage_inst_dmem_ram_213__0_), .D(
        mem_stage_inst_dmem_ram_215__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n239) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1240 ( .A(
        mem_stage_inst_dmem_ram_220__0_), .B(mem_stage_inst_dmem_ram_222__0_), 
        .C(mem_stage_inst_dmem_ram_221__0_), .D(
        mem_stage_inst_dmem_ram_223__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n240) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1239 ( .A(mem_stage_inst_dmem_n237), 
        .B(mem_stage_inst_dmem_n238), .C(mem_stage_inst_dmem_n239), .D(
        mem_stage_inst_dmem_n240), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n236) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1238 ( .A(
        mem_stage_inst_dmem_ram_80__0_), .B(mem_stage_inst_dmem_ram_82__0_), 
        .C(mem_stage_inst_dmem_ram_81__0_), .D(mem_stage_inst_dmem_ram_83__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n277) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1237 ( .A(
        mem_stage_inst_dmem_ram_84__0_), .B(mem_stage_inst_dmem_ram_86__0_), 
        .C(mem_stage_inst_dmem_ram_85__0_), .D(mem_stage_inst_dmem_ram_87__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n279) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1236 ( .A(
        mem_stage_inst_dmem_ram_92__0_), .B(mem_stage_inst_dmem_ram_94__0_), 
        .C(mem_stage_inst_dmem_ram_93__0_), .D(mem_stage_inst_dmem_ram_95__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n280) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1235 ( .A(mem_stage_inst_dmem_n277), 
        .B(mem_stage_inst_dmem_n278), .C(mem_stage_inst_dmem_n279), .D(
        mem_stage_inst_dmem_n280), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n276) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1234 ( .A(
        mem_stage_inst_dmem_ram_52__15_), .B(mem_stage_inst_dmem_ram_54__15_), 
        .C(mem_stage_inst_dmem_ram_53__15_), .D(
        mem_stage_inst_dmem_ram_55__15_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n2), .Y(mem_stage_inst_dmem_n5645) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1233 ( .A(
        mem_stage_inst_dmem_ram_20__15_), .B(mem_stage_inst_dmem_ram_22__15_), 
        .C(mem_stage_inst_dmem_ram_21__15_), .D(
        mem_stage_inst_dmem_ram_23__15_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n5655) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1232 ( .A(
        mem_stage_inst_dmem_ram_4__15_), .B(mem_stage_inst_dmem_ram_6__15_), 
        .C(mem_stage_inst_dmem_ram_5__15_), .D(mem_stage_inst_dmem_ram_7__15_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n5660) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1231 ( .A(
        mem_stage_inst_dmem_ram_180__15_), .B(mem_stage_inst_dmem_ram_182__15_), .C(mem_stage_inst_dmem_ram_181__15_), .D(mem_stage_inst_dmem_ram_183__15_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5605) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1230 ( .A(
        mem_stage_inst_dmem_ram_148__15_), .B(mem_stage_inst_dmem_ram_150__15_), .C(mem_stage_inst_dmem_ram_149__15_), .D(mem_stage_inst_dmem_ram_151__15_), 
        .S0(mem_stage_inst_dmem_n154), .S1(mem_stage_inst_dmem_n4), .Y(
        mem_stage_inst_dmem_n5615) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1229 ( .A(
        mem_stage_inst_dmem_ram_132__15_), .B(mem_stage_inst_dmem_ram_134__15_), .C(mem_stage_inst_dmem_ram_133__15_), .D(mem_stage_inst_dmem_ram_135__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5620) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1228 ( .A(
        mem_stage_inst_dmem_ram_52__14_), .B(mem_stage_inst_dmem_ram_54__14_), 
        .C(mem_stage_inst_dmem_ram_53__14_), .D(
        mem_stage_inst_dmem_ram_55__14_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5561) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1227 ( .A(
        mem_stage_inst_dmem_ram_20__14_), .B(mem_stage_inst_dmem_ram_22__14_), 
        .C(mem_stage_inst_dmem_ram_21__14_), .D(
        mem_stage_inst_dmem_ram_23__14_), .S0(mem_stage_inst_dmem_n101), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5571) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1226 ( .A(
        mem_stage_inst_dmem_ram_4__14_), .B(mem_stage_inst_dmem_ram_6__14_), 
        .C(mem_stage_inst_dmem_ram_5__14_), .D(mem_stage_inst_dmem_ram_7__14_), 
        .S0(mem_stage_inst_dmem_n102), .S1(mem_stage_inst_dmem_n27), .Y(
        mem_stage_inst_dmem_n5576) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1225 ( .A(
        mem_stage_inst_dmem_ram_180__14_), .B(mem_stage_inst_dmem_ram_182__14_), .C(mem_stage_inst_dmem_ram_181__14_), .D(mem_stage_inst_dmem_ram_183__14_), 
        .S0(mem_stage_inst_dmem_n114), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5521) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1224 ( .A(
        mem_stage_inst_dmem_ram_148__14_), .B(mem_stage_inst_dmem_ram_150__14_), .C(mem_stage_inst_dmem_ram_149__14_), .D(mem_stage_inst_dmem_ram_151__14_), 
        .S0(mem_stage_inst_dmem_n115), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5531) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1223 ( .A(
        mem_stage_inst_dmem_ram_132__14_), .B(mem_stage_inst_dmem_ram_134__14_), .C(mem_stage_inst_dmem_ram_133__14_), .D(mem_stage_inst_dmem_ram_135__14_), 
        .S0(mem_stage_inst_dmem_n150), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5536) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1222 ( .A(
        mem_stage_inst_dmem_ram_52__13_), .B(mem_stage_inst_dmem_ram_54__13_), 
        .C(mem_stage_inst_dmem_ram_53__13_), .D(
        mem_stage_inst_dmem_ram_55__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5477) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1221 ( .A(
        mem_stage_inst_dmem_ram_20__13_), .B(mem_stage_inst_dmem_ram_22__13_), 
        .C(mem_stage_inst_dmem_ram_21__13_), .D(
        mem_stage_inst_dmem_ram_23__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5487) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1220 ( .A(
        mem_stage_inst_dmem_ram_4__13_), .B(mem_stage_inst_dmem_ram_6__13_), 
        .C(mem_stage_inst_dmem_ram_5__13_), .D(mem_stage_inst_dmem_ram_7__13_), 
        .S0(mem_stage_inst_dmem_n125), .S1(mem_stage_inst_dmem_n27), .Y(
        mem_stage_inst_dmem_n5492) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1219 ( .A(
        mem_stage_inst_dmem_ram_180__13_), .B(mem_stage_inst_dmem_ram_182__13_), .C(mem_stage_inst_dmem_ram_181__13_), .D(mem_stage_inst_dmem_ram_183__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n34), .Y(
        mem_stage_inst_dmem_n5437) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1218 ( .A(
        mem_stage_inst_dmem_ram_148__13_), .B(mem_stage_inst_dmem_ram_150__13_), .C(mem_stage_inst_dmem_ram_149__13_), .D(mem_stage_inst_dmem_ram_151__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5447) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1217 ( .A(
        mem_stage_inst_dmem_ram_132__13_), .B(mem_stage_inst_dmem_ram_134__13_), .C(mem_stage_inst_dmem_ram_133__13_), .D(mem_stage_inst_dmem_ram_135__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5452) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1216 ( .A(
        mem_stage_inst_dmem_ram_52__12_), .B(mem_stage_inst_dmem_ram_54__12_), 
        .C(mem_stage_inst_dmem_ram_53__12_), .D(
        mem_stage_inst_dmem_ram_55__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n5393) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1215 ( .A(
        mem_stage_inst_dmem_ram_20__12_), .B(mem_stage_inst_dmem_ram_22__12_), 
        .C(mem_stage_inst_dmem_ram_21__12_), .D(
        mem_stage_inst_dmem_ram_23__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n5403) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1214 ( .A(
        mem_stage_inst_dmem_ram_4__12_), .B(mem_stage_inst_dmem_ram_6__12_), 
        .C(mem_stage_inst_dmem_ram_5__12_), .D(mem_stage_inst_dmem_ram_7__12_), 
        .S0(mem_stage_inst_dmem_n141), .S1(mem_stage_inst_dmem_n13), .Y(
        mem_stage_inst_dmem_n5408) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1213 ( .A(
        mem_stage_inst_dmem_ram_180__12_), .B(mem_stage_inst_dmem_ram_182__12_), .C(mem_stage_inst_dmem_ram_181__12_), .D(mem_stage_inst_dmem_ram_183__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5353) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1212 ( .A(
        mem_stage_inst_dmem_ram_148__12_), .B(mem_stage_inst_dmem_ram_150__12_), .C(mem_stage_inst_dmem_ram_149__12_), .D(mem_stage_inst_dmem_ram_151__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5363) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1211 ( .A(
        mem_stage_inst_dmem_ram_132__12_), .B(mem_stage_inst_dmem_ram_134__12_), .C(mem_stage_inst_dmem_ram_133__12_), .D(mem_stage_inst_dmem_ram_135__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5368) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1210 ( .A(
        mem_stage_inst_dmem_ram_52__11_), .B(mem_stage_inst_dmem_ram_54__11_), 
        .C(mem_stage_inst_dmem_ram_53__11_), .D(
        mem_stage_inst_dmem_ram_55__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5309) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1209 ( .A(
        mem_stage_inst_dmem_ram_20__11_), .B(mem_stage_inst_dmem_ram_22__11_), 
        .C(mem_stage_inst_dmem_ram_21__11_), .D(
        mem_stage_inst_dmem_ram_23__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5319) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1208 ( .A(
        mem_stage_inst_dmem_ram_4__11_), .B(mem_stage_inst_dmem_ram_6__11_), 
        .C(mem_stage_inst_dmem_ram_5__11_), .D(mem_stage_inst_dmem_ram_7__11_), 
        .S0(mem_stage_inst_dmem_n108), .S1(mem_stage_inst_dmem_n10), .Y(
        mem_stage_inst_dmem_n5324) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1207 ( .A(
        mem_stage_inst_dmem_ram_180__11_), .B(mem_stage_inst_dmem_ram_182__11_), .C(mem_stage_inst_dmem_ram_181__11_), .D(mem_stage_inst_dmem_ram_183__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5269) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1206 ( .A(
        mem_stage_inst_dmem_ram_148__11_), .B(mem_stage_inst_dmem_ram_150__11_), .C(mem_stage_inst_dmem_ram_149__11_), .D(mem_stage_inst_dmem_ram_151__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5279) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1205 ( .A(
        mem_stage_inst_dmem_ram_132__11_), .B(mem_stage_inst_dmem_ram_134__11_), .C(mem_stage_inst_dmem_ram_133__11_), .D(mem_stage_inst_dmem_ram_135__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5284) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1204 ( .A(
        mem_stage_inst_dmem_ram_52__10_), .B(mem_stage_inst_dmem_ram_54__10_), 
        .C(mem_stage_inst_dmem_ram_53__10_), .D(
        mem_stage_inst_dmem_ram_55__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5225) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1203 ( .A(
        mem_stage_inst_dmem_ram_20__10_), .B(mem_stage_inst_dmem_ram_22__10_), 
        .C(mem_stage_inst_dmem_ram_21__10_), .D(
        mem_stage_inst_dmem_ram_23__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5235) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1202 ( .A(
        mem_stage_inst_dmem_ram_4__10_), .B(mem_stage_inst_dmem_ram_6__10_), 
        .C(mem_stage_inst_dmem_ram_5__10_), .D(mem_stage_inst_dmem_ram_7__10_), 
        .S0(mem_stage_inst_dmem_n103), .S1(mem_stage_inst_dmem_n5), .Y(
        mem_stage_inst_dmem_n5240) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1201 ( .A(
        mem_stage_inst_dmem_ram_180__10_), .B(mem_stage_inst_dmem_ram_182__10_), .C(mem_stage_inst_dmem_ram_181__10_), .D(mem_stage_inst_dmem_ram_183__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5185) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1200 ( .A(
        mem_stage_inst_dmem_ram_148__10_), .B(mem_stage_inst_dmem_ram_150__10_), .C(mem_stage_inst_dmem_ram_149__10_), .D(mem_stage_inst_dmem_ram_151__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5195) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1199 ( .A(
        mem_stage_inst_dmem_ram_132__10_), .B(mem_stage_inst_dmem_ram_134__10_), .C(mem_stage_inst_dmem_ram_133__10_), .D(mem_stage_inst_dmem_ram_135__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5200) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1198 ( .A(
        mem_stage_inst_dmem_ram_52__9_), .B(mem_stage_inst_dmem_ram_54__9_), 
        .C(mem_stage_inst_dmem_ram_53__9_), .D(mem_stage_inst_dmem_ram_55__9_), 
        .S0(mem_stage_inst_dmem_n139), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n5141) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1197 ( .A(
        mem_stage_inst_dmem_ram_20__9_), .B(mem_stage_inst_dmem_ram_22__9_), 
        .C(mem_stage_inst_dmem_ram_21__9_), .D(mem_stage_inst_dmem_ram_23__9_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n43), .Y(
        mem_stage_inst_dmem_n5151) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1196 ( .A(mem_stage_inst_dmem_ram_4__9_), .B(mem_stage_inst_dmem_ram_6__9_), .C(mem_stage_inst_dmem_ram_5__9_), .D(
        mem_stage_inst_dmem_ram_7__9_), .S0(mem_stage_inst_dmem_n164), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n5156) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1195 ( .A(
        mem_stage_inst_dmem_ram_180__9_), .B(mem_stage_inst_dmem_ram_182__9_), 
        .C(mem_stage_inst_dmem_ram_181__9_), .D(
        mem_stage_inst_dmem_ram_183__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5101) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1194 ( .A(
        mem_stage_inst_dmem_ram_148__9_), .B(mem_stage_inst_dmem_ram_150__9_), 
        .C(mem_stage_inst_dmem_ram_149__9_), .D(
        mem_stage_inst_dmem_ram_151__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5111) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1193 ( .A(
        mem_stage_inst_dmem_ram_132__9_), .B(mem_stage_inst_dmem_ram_134__9_), 
        .C(mem_stage_inst_dmem_ram_133__9_), .D(
        mem_stage_inst_dmem_ram_135__9_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5116) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1192 ( .A(
        mem_stage_inst_dmem_ram_52__8_), .B(mem_stage_inst_dmem_ram_54__8_), 
        .C(mem_stage_inst_dmem_ram_53__8_), .D(mem_stage_inst_dmem_ram_55__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5057) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1191 ( .A(
        mem_stage_inst_dmem_ram_20__8_), .B(mem_stage_inst_dmem_ram_22__8_), 
        .C(mem_stage_inst_dmem_ram_21__8_), .D(mem_stage_inst_dmem_ram_23__8_), 
        .S0(mem_stage_inst_dmem_n113), .S1(mem_stage_inst_dmem_n15), .Y(
        mem_stage_inst_dmem_n5067) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1190 ( .A(mem_stage_inst_dmem_ram_4__8_), .B(mem_stage_inst_dmem_ram_6__8_), .C(mem_stage_inst_dmem_ram_5__8_), .D(
        mem_stage_inst_dmem_ram_7__8_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5072) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1189 ( .A(
        mem_stage_inst_dmem_ram_180__8_), .B(mem_stage_inst_dmem_ram_182__8_), 
        .C(mem_stage_inst_dmem_ram_181__8_), .D(
        mem_stage_inst_dmem_ram_183__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5017) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1188 ( .A(
        mem_stage_inst_dmem_ram_148__8_), .B(mem_stage_inst_dmem_ram_150__8_), 
        .C(mem_stage_inst_dmem_ram_149__8_), .D(
        mem_stage_inst_dmem_ram_151__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5027) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1187 ( .A(
        mem_stage_inst_dmem_ram_132__8_), .B(mem_stage_inst_dmem_ram_134__8_), 
        .C(mem_stage_inst_dmem_ram_133__8_), .D(
        mem_stage_inst_dmem_ram_135__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5032) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1186 ( .A(
        mem_stage_inst_dmem_ram_52__7_), .B(mem_stage_inst_dmem_ram_54__7_), 
        .C(mem_stage_inst_dmem_ram_53__7_), .D(mem_stage_inst_dmem_ram_55__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4973) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1185 ( .A(
        mem_stage_inst_dmem_ram_20__7_), .B(mem_stage_inst_dmem_ram_22__7_), 
        .C(mem_stage_inst_dmem_ram_21__7_), .D(mem_stage_inst_dmem_ram_23__7_), 
        .S0(mem_stage_inst_dmem_n154), .S1(mem_stage_inst_dmem_n56), .Y(
        mem_stage_inst_dmem_n4983) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1184 ( .A(mem_stage_inst_dmem_ram_4__7_), .B(mem_stage_inst_dmem_ram_6__7_), .C(mem_stage_inst_dmem_ram_5__7_), .D(
        mem_stage_inst_dmem_ram_7__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4988) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1183 ( .A(
        mem_stage_inst_dmem_ram_180__7_), .B(mem_stage_inst_dmem_ram_182__7_), 
        .C(mem_stage_inst_dmem_ram_181__7_), .D(
        mem_stage_inst_dmem_ram_183__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4933) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1182 ( .A(
        mem_stage_inst_dmem_ram_148__7_), .B(mem_stage_inst_dmem_ram_150__7_), 
        .C(mem_stage_inst_dmem_ram_149__7_), .D(
        mem_stage_inst_dmem_ram_151__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4943) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1181 ( .A(
        mem_stage_inst_dmem_ram_132__7_), .B(mem_stage_inst_dmem_ram_134__7_), 
        .C(mem_stage_inst_dmem_ram_133__7_), .D(
        mem_stage_inst_dmem_ram_135__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4948) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1180 ( .A(
        mem_stage_inst_dmem_ram_52__6_), .B(mem_stage_inst_dmem_ram_54__6_), 
        .C(mem_stage_inst_dmem_ram_53__6_), .D(mem_stage_inst_dmem_ram_55__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4889) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1179 ( .A(
        mem_stage_inst_dmem_ram_20__6_), .B(mem_stage_inst_dmem_ram_22__6_), 
        .C(mem_stage_inst_dmem_ram_21__6_), .D(mem_stage_inst_dmem_ram_23__6_), 
        .S0(mem_stage_inst_dmem_n149), .S1(mem_stage_inst_dmem_n51), .Y(
        mem_stage_inst_dmem_n4899) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1178 ( .A(mem_stage_inst_dmem_ram_4__6_), .B(mem_stage_inst_dmem_ram_6__6_), .C(mem_stage_inst_dmem_ram_5__6_), .D(
        mem_stage_inst_dmem_ram_7__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4904) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1177 ( .A(
        mem_stage_inst_dmem_ram_180__6_), .B(mem_stage_inst_dmem_ram_182__6_), 
        .C(mem_stage_inst_dmem_ram_181__6_), .D(
        mem_stage_inst_dmem_ram_183__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4849) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1176 ( .A(
        mem_stage_inst_dmem_ram_148__6_), .B(mem_stage_inst_dmem_ram_150__6_), 
        .C(mem_stage_inst_dmem_ram_149__6_), .D(
        mem_stage_inst_dmem_ram_151__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4859) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1175 ( .A(
        mem_stage_inst_dmem_ram_132__6_), .B(mem_stage_inst_dmem_ram_134__6_), 
        .C(mem_stage_inst_dmem_ram_133__6_), .D(
        mem_stage_inst_dmem_ram_135__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4864) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1174 ( .A(
        mem_stage_inst_dmem_ram_52__5_), .B(mem_stage_inst_dmem_ram_54__5_), 
        .C(mem_stage_inst_dmem_ram_53__5_), .D(mem_stage_inst_dmem_ram_55__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4805) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1173 ( .A(
        mem_stage_inst_dmem_ram_20__5_), .B(mem_stage_inst_dmem_ram_22__5_), 
        .C(mem_stage_inst_dmem_ram_21__5_), .D(mem_stage_inst_dmem_ram_23__5_), 
        .S0(mem_stage_inst_dmem_n164), .S1(ex_pipeline_reg_out[22]), .Y(
        mem_stage_inst_dmem_n4815) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1172 ( .A(mem_stage_inst_dmem_ram_4__5_), .B(mem_stage_inst_dmem_ram_6__5_), .C(mem_stage_inst_dmem_ram_5__5_), .D(
        mem_stage_inst_dmem_ram_7__5_), .S0(mem_stage_inst_dmem_n164), .S1(
        ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4820) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1171 ( .A(
        mem_stage_inst_dmem_ram_180__5_), .B(mem_stage_inst_dmem_ram_182__5_), 
        .C(mem_stage_inst_dmem_ram_181__5_), .D(
        mem_stage_inst_dmem_ram_183__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4765) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1170 ( .A(
        mem_stage_inst_dmem_ram_148__5_), .B(mem_stage_inst_dmem_ram_150__5_), 
        .C(mem_stage_inst_dmem_ram_149__5_), .D(
        mem_stage_inst_dmem_ram_151__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4775) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1169 ( .A(
        mem_stage_inst_dmem_ram_132__5_), .B(mem_stage_inst_dmem_ram_134__5_), 
        .C(mem_stage_inst_dmem_ram_133__5_), .D(
        mem_stage_inst_dmem_ram_135__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4780) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1168 ( .A(
        mem_stage_inst_dmem_ram_52__4_), .B(mem_stage_inst_dmem_ram_54__4_), 
        .C(mem_stage_inst_dmem_ram_53__4_), .D(mem_stage_inst_dmem_ram_55__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4721) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1167 ( .A(
        mem_stage_inst_dmem_ram_20__4_), .B(mem_stage_inst_dmem_ram_22__4_), 
        .C(mem_stage_inst_dmem_ram_21__4_), .D(mem_stage_inst_dmem_ram_23__4_), 
        .S0(mem_stage_inst_dmem_n159), .S1(mem_stage_inst_dmem_n61), .Y(
        mem_stage_inst_dmem_n4731) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1166 ( .A(mem_stage_inst_dmem_ram_4__4_), .B(mem_stage_inst_dmem_ram_6__4_), .C(mem_stage_inst_dmem_ram_5__4_), .D(
        mem_stage_inst_dmem_ram_7__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4736) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1165 ( .A(
        mem_stage_inst_dmem_ram_180__4_), .B(mem_stage_inst_dmem_ram_182__4_), 
        .C(mem_stage_inst_dmem_ram_181__4_), .D(
        mem_stage_inst_dmem_ram_183__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4681) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1164 ( .A(
        mem_stage_inst_dmem_ram_148__4_), .B(mem_stage_inst_dmem_ram_150__4_), 
        .C(mem_stage_inst_dmem_ram_149__4_), .D(
        mem_stage_inst_dmem_ram_151__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4691) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1163 ( .A(
        mem_stage_inst_dmem_ram_132__4_), .B(mem_stage_inst_dmem_ram_134__4_), 
        .C(mem_stage_inst_dmem_ram_133__4_), .D(
        mem_stage_inst_dmem_ram_135__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4696) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1162 ( .A(
        mem_stage_inst_dmem_ram_52__3_), .B(mem_stage_inst_dmem_ram_54__3_), 
        .C(mem_stage_inst_dmem_ram_53__3_), .D(mem_stage_inst_dmem_ram_55__3_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n541) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1161 ( .A(
        mem_stage_inst_dmem_ram_20__3_), .B(mem_stage_inst_dmem_ram_22__3_), 
        .C(mem_stage_inst_dmem_ram_21__3_), .D(mem_stage_inst_dmem_ram_23__3_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n551) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1160 ( .A(mem_stage_inst_dmem_ram_4__3_), .B(mem_stage_inst_dmem_ram_6__3_), .C(mem_stage_inst_dmem_ram_5__3_), .D(
        mem_stage_inst_dmem_ram_7__3_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n556) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1159 ( .A(
        mem_stage_inst_dmem_ram_180__3_), .B(mem_stage_inst_dmem_ram_182__3_), 
        .C(mem_stage_inst_dmem_ram_181__3_), .D(
        mem_stage_inst_dmem_ram_183__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n501) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1158 ( .A(
        mem_stage_inst_dmem_ram_148__3_), .B(mem_stage_inst_dmem_ram_150__3_), 
        .C(mem_stage_inst_dmem_ram_149__3_), .D(
        mem_stage_inst_dmem_ram_151__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n511) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1157 ( .A(
        mem_stage_inst_dmem_ram_132__3_), .B(mem_stage_inst_dmem_ram_134__3_), 
        .C(mem_stage_inst_dmem_ram_133__3_), .D(
        mem_stage_inst_dmem_ram_135__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n516) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1156 ( .A(
        mem_stage_inst_dmem_ram_52__2_), .B(mem_stage_inst_dmem_ram_54__2_), 
        .C(mem_stage_inst_dmem_ram_53__2_), .D(mem_stage_inst_dmem_ram_55__2_), 
        .S0(mem_stage_inst_dmem_n129), .S1(mem_stage_inst_dmem_n31), .Y(
        mem_stage_inst_dmem_n457) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1155 ( .A(
        mem_stage_inst_dmem_ram_20__2_), .B(mem_stage_inst_dmem_ram_22__2_), 
        .C(mem_stage_inst_dmem_ram_21__2_), .D(mem_stage_inst_dmem_ram_23__2_), 
        .S0(mem_stage_inst_dmem_n129), .S1(mem_stage_inst_dmem_n31), .Y(
        mem_stage_inst_dmem_n467) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1154 ( .A(mem_stage_inst_dmem_ram_4__2_), .B(mem_stage_inst_dmem_ram_6__2_), .C(mem_stage_inst_dmem_ram_5__2_), .D(
        mem_stage_inst_dmem_ram_7__2_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n472) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1153 ( .A(
        mem_stage_inst_dmem_ram_180__2_), .B(mem_stage_inst_dmem_ram_182__2_), 
        .C(mem_stage_inst_dmem_ram_181__2_), .D(
        mem_stage_inst_dmem_ram_183__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n417) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1152 ( .A(
        mem_stage_inst_dmem_ram_148__2_), .B(mem_stage_inst_dmem_ram_150__2_), 
        .C(mem_stage_inst_dmem_ram_149__2_), .D(
        mem_stage_inst_dmem_ram_151__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n427) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1151 ( .A(
        mem_stage_inst_dmem_ram_132__2_), .B(mem_stage_inst_dmem_ram_134__2_), 
        .C(mem_stage_inst_dmem_ram_133__2_), .D(
        mem_stage_inst_dmem_ram_135__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n432) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1150 ( .A(
        mem_stage_inst_dmem_ram_52__1_), .B(mem_stage_inst_dmem_ram_54__1_), 
        .C(mem_stage_inst_dmem_ram_53__1_), .D(mem_stage_inst_dmem_ram_55__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n373) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1149 ( .A(
        mem_stage_inst_dmem_ram_20__1_), .B(mem_stage_inst_dmem_ram_22__1_), 
        .C(mem_stage_inst_dmem_ram_21__1_), .D(mem_stage_inst_dmem_ram_23__1_), 
        .S0(mem_stage_inst_dmem_n144), .S1(mem_stage_inst_dmem_n46), .Y(
        mem_stage_inst_dmem_n383) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1148 ( .A(mem_stage_inst_dmem_ram_4__1_), .B(mem_stage_inst_dmem_ram_6__1_), .C(mem_stage_inst_dmem_ram_5__1_), .D(
        mem_stage_inst_dmem_ram_7__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n388) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1147 ( .A(
        mem_stage_inst_dmem_ram_180__1_), .B(mem_stage_inst_dmem_ram_182__1_), 
        .C(mem_stage_inst_dmem_ram_181__1_), .D(
        mem_stage_inst_dmem_ram_183__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n333) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1146 ( .A(
        mem_stage_inst_dmem_ram_148__1_), .B(mem_stage_inst_dmem_ram_150__1_), 
        .C(mem_stage_inst_dmem_ram_149__1_), .D(
        mem_stage_inst_dmem_ram_151__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n343) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1145 ( .A(
        mem_stage_inst_dmem_ram_132__1_), .B(mem_stage_inst_dmem_ram_134__1_), 
        .C(mem_stage_inst_dmem_ram_133__1_), .D(
        mem_stage_inst_dmem_ram_135__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n348) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1144 ( .A(
        mem_stage_inst_dmem_ram_52__0_), .B(mem_stage_inst_dmem_ram_54__0_), 
        .C(mem_stage_inst_dmem_ram_53__0_), .D(mem_stage_inst_dmem_ram_55__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n289) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1143 ( .A(
        mem_stage_inst_dmem_ram_20__0_), .B(mem_stage_inst_dmem_ram_22__0_), 
        .C(mem_stage_inst_dmem_ram_21__0_), .D(mem_stage_inst_dmem_ram_23__0_), 
        .S0(mem_stage_inst_dmem_n139), .S1(mem_stage_inst_dmem_n41), .Y(
        mem_stage_inst_dmem_n299) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1142 ( .A(mem_stage_inst_dmem_ram_4__0_), .B(mem_stage_inst_dmem_ram_6__0_), .C(mem_stage_inst_dmem_ram_5__0_), .D(
        mem_stage_inst_dmem_ram_7__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n304) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1141 ( .A(
        mem_stage_inst_dmem_ram_180__0_), .B(mem_stage_inst_dmem_ram_182__0_), 
        .C(mem_stage_inst_dmem_ram_181__0_), .D(
        mem_stage_inst_dmem_ram_183__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n249) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1140 ( .A(
        mem_stage_inst_dmem_ram_148__0_), .B(mem_stage_inst_dmem_ram_150__0_), 
        .C(mem_stage_inst_dmem_ram_149__0_), .D(
        mem_stage_inst_dmem_ram_151__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n259) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1139 ( .A(
        mem_stage_inst_dmem_ram_132__0_), .B(mem_stage_inst_dmem_ram_134__0_), 
        .C(mem_stage_inst_dmem_ram_133__0_), .D(
        mem_stage_inst_dmem_ram_135__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n264) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1138 ( .A(
        mem_stage_inst_dmem_ram_192__15_), .B(mem_stage_inst_dmem_ram_194__15_), .C(mem_stage_inst_dmem_ram_193__15_), .D(mem_stage_inst_dmem_ram_195__15_), 
        .S0(mem_stage_inst_dmem_n132), .S1(mem_stage_inst_dmem_n15), .Y(
        mem_stage_inst_dmem_n5598) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1137 ( .A(
        mem_stage_inst_dmem_ram_196__15_), .B(mem_stage_inst_dmem_ram_198__15_), .C(mem_stage_inst_dmem_ram_197__15_), .D(mem_stage_inst_dmem_ram_199__15_), 
        .S0(mem_stage_inst_dmem_n131), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5600) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1136 ( .A(
        mem_stage_inst_dmem_ram_204__15_), .B(mem_stage_inst_dmem_ram_206__15_), .C(mem_stage_inst_dmem_ram_205__15_), .D(mem_stage_inst_dmem_ram_207__15_), 
        .S0(mem_stage_inst_dmem_n130), .S1(mem_stage_inst_dmem_n41), .Y(
        mem_stage_inst_dmem_n5601) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1135 ( .A(mem_stage_inst_dmem_n5598), 
        .B(mem_stage_inst_dmem_n5599), .C(mem_stage_inst_dmem_n5600), .D(
        mem_stage_inst_dmem_n5601), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5597) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1134 ( .A(
        mem_stage_inst_dmem_ram_64__15_), .B(mem_stage_inst_dmem_ram_66__15_), 
        .C(mem_stage_inst_dmem_ram_65__15_), .D(
        mem_stage_inst_dmem_ram_67__15_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n5638) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1133 ( .A(
        mem_stage_inst_dmem_ram_68__15_), .B(mem_stage_inst_dmem_ram_70__15_), 
        .C(mem_stage_inst_dmem_ram_69__15_), .D(
        mem_stage_inst_dmem_ram_71__15_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n5640) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1132 ( .A(
        mem_stage_inst_dmem_ram_76__15_), .B(mem_stage_inst_dmem_ram_78__15_), 
        .C(mem_stage_inst_dmem_ram_77__15_), .D(
        mem_stage_inst_dmem_ram_79__15_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n5641) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1131 ( .A(mem_stage_inst_dmem_n5638), 
        .B(mem_stage_inst_dmem_n5639), .C(mem_stage_inst_dmem_n5640), .D(
        mem_stage_inst_dmem_n5641), .S0(mem_stage_inst_dmem_n212), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5637) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1130 ( .A(
        mem_stage_inst_dmem_ram_192__14_), .B(mem_stage_inst_dmem_ram_194__14_), .C(mem_stage_inst_dmem_ram_193__14_), .D(mem_stage_inst_dmem_ram_195__14_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n53), .Y(
        mem_stage_inst_dmem_n5514) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1129 ( .A(
        mem_stage_inst_dmem_ram_196__14_), .B(mem_stage_inst_dmem_ram_198__14_), .C(mem_stage_inst_dmem_ram_197__14_), .D(mem_stage_inst_dmem_ram_199__14_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n52), .Y(
        mem_stage_inst_dmem_n5516) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1128 ( .A(
        mem_stage_inst_dmem_ram_204__14_), .B(mem_stage_inst_dmem_ram_206__14_), .C(mem_stage_inst_dmem_ram_205__14_), .D(mem_stage_inst_dmem_ram_207__14_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n39), .Y(
        mem_stage_inst_dmem_n5517) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1127 ( .A(mem_stage_inst_dmem_n5514), 
        .B(mem_stage_inst_dmem_n5515), .C(mem_stage_inst_dmem_n5516), .D(
        mem_stage_inst_dmem_n5517), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5513) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1126 ( .A(
        mem_stage_inst_dmem_ram_64__14_), .B(mem_stage_inst_dmem_ram_66__14_), 
        .C(mem_stage_inst_dmem_ram_65__14_), .D(
        mem_stage_inst_dmem_ram_67__14_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5554) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1125 ( .A(
        mem_stage_inst_dmem_ram_68__14_), .B(mem_stage_inst_dmem_ram_70__14_), 
        .C(mem_stage_inst_dmem_ram_69__14_), .D(
        mem_stage_inst_dmem_ram_71__14_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5556) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1124 ( .A(
        mem_stage_inst_dmem_ram_76__14_), .B(mem_stage_inst_dmem_ram_78__14_), 
        .C(mem_stage_inst_dmem_ram_77__14_), .D(
        mem_stage_inst_dmem_ram_79__14_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5557) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1123 ( .A(mem_stage_inst_dmem_n5554), 
        .B(mem_stage_inst_dmem_n5555), .C(mem_stage_inst_dmem_n5556), .D(
        mem_stage_inst_dmem_n5557), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5553) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1122 ( .A(
        mem_stage_inst_dmem_ram_192__13_), .B(mem_stage_inst_dmem_ram_194__13_), .C(mem_stage_inst_dmem_ram_193__13_), .D(mem_stage_inst_dmem_ram_195__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n5430) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1121 ( .A(
        mem_stage_inst_dmem_ram_196__13_), .B(mem_stage_inst_dmem_ram_198__13_), .C(mem_stage_inst_dmem_ram_197__13_), .D(mem_stage_inst_dmem_ram_199__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n39), .Y(
        mem_stage_inst_dmem_n5432) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1120 ( .A(
        mem_stage_inst_dmem_ram_204__13_), .B(mem_stage_inst_dmem_ram_206__13_), .C(mem_stage_inst_dmem_ram_205__13_), .D(mem_stage_inst_dmem_ram_207__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n38), .Y(
        mem_stage_inst_dmem_n5433) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1119 ( .A(mem_stage_inst_dmem_n5430), 
        .B(mem_stage_inst_dmem_n5431), .C(mem_stage_inst_dmem_n5432), .D(
        mem_stage_inst_dmem_n5433), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5429) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1118 ( .A(
        mem_stage_inst_dmem_ram_64__13_), .B(mem_stage_inst_dmem_ram_66__13_), 
        .C(mem_stage_inst_dmem_ram_65__13_), .D(
        mem_stage_inst_dmem_ram_67__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5470) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1117 ( .A(
        mem_stage_inst_dmem_ram_68__13_), .B(mem_stage_inst_dmem_ram_70__13_), 
        .C(mem_stage_inst_dmem_ram_69__13_), .D(
        mem_stage_inst_dmem_ram_71__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5472) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1116 ( .A(
        mem_stage_inst_dmem_ram_76__13_), .B(mem_stage_inst_dmem_ram_78__13_), 
        .C(mem_stage_inst_dmem_ram_77__13_), .D(
        mem_stage_inst_dmem_ram_79__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n5473) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1115 ( .A(mem_stage_inst_dmem_n5470), 
        .B(mem_stage_inst_dmem_n5471), .C(mem_stage_inst_dmem_n5472), .D(
        mem_stage_inst_dmem_n5473), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5469) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1114 ( .A(
        mem_stage_inst_dmem_ram_192__12_), .B(mem_stage_inst_dmem_ram_194__12_), .C(mem_stage_inst_dmem_ram_193__12_), .D(mem_stage_inst_dmem_ram_195__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5346) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1113 ( .A(
        mem_stage_inst_dmem_ram_196__12_), .B(mem_stage_inst_dmem_ram_198__12_), .C(mem_stage_inst_dmem_ram_197__12_), .D(mem_stage_inst_dmem_ram_199__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5348) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1112 ( .A(
        mem_stage_inst_dmem_ram_204__12_), .B(mem_stage_inst_dmem_ram_206__12_), .C(mem_stage_inst_dmem_ram_205__12_), .D(mem_stage_inst_dmem_ram_207__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5349) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1111 ( .A(mem_stage_inst_dmem_n5346), 
        .B(mem_stage_inst_dmem_n5347), .C(mem_stage_inst_dmem_n5348), .D(
        mem_stage_inst_dmem_n5349), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5345) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1110 ( .A(
        mem_stage_inst_dmem_ram_64__12_), .B(mem_stage_inst_dmem_ram_66__12_), 
        .C(mem_stage_inst_dmem_ram_65__12_), .D(
        mem_stage_inst_dmem_ram_67__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n5386) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1109 ( .A(
        mem_stage_inst_dmem_ram_68__12_), .B(mem_stage_inst_dmem_ram_70__12_), 
        .C(mem_stage_inst_dmem_ram_69__12_), .D(
        mem_stage_inst_dmem_ram_71__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n5388) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1108 ( .A(
        mem_stage_inst_dmem_ram_76__12_), .B(mem_stage_inst_dmem_ram_78__12_), 
        .C(mem_stage_inst_dmem_ram_77__12_), .D(
        mem_stage_inst_dmem_ram_79__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5389) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1107 ( .A(mem_stage_inst_dmem_n5386), 
        .B(mem_stage_inst_dmem_n5387), .C(mem_stage_inst_dmem_n5388), .D(
        mem_stage_inst_dmem_n5389), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5385) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1106 ( .A(
        mem_stage_inst_dmem_ram_192__11_), .B(mem_stage_inst_dmem_ram_194__11_), .C(mem_stage_inst_dmem_ram_193__11_), .D(mem_stage_inst_dmem_ram_195__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5262) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1105 ( .A(
        mem_stage_inst_dmem_ram_196__11_), .B(mem_stage_inst_dmem_ram_198__11_), .C(mem_stage_inst_dmem_ram_197__11_), .D(mem_stage_inst_dmem_ram_199__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5264) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1104 ( .A(
        mem_stage_inst_dmem_ram_204__11_), .B(mem_stage_inst_dmem_ram_206__11_), .C(mem_stage_inst_dmem_ram_205__11_), .D(mem_stage_inst_dmem_ram_207__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5265) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1103 ( .A(mem_stage_inst_dmem_n5262), 
        .B(mem_stage_inst_dmem_n5263), .C(mem_stage_inst_dmem_n5264), .D(
        mem_stage_inst_dmem_n5265), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5261) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1102 ( .A(
        mem_stage_inst_dmem_ram_64__11_), .B(mem_stage_inst_dmem_ram_66__11_), 
        .C(mem_stage_inst_dmem_ram_65__11_), .D(
        mem_stage_inst_dmem_ram_67__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5302) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1101 ( .A(
        mem_stage_inst_dmem_ram_68__11_), .B(mem_stage_inst_dmem_ram_70__11_), 
        .C(mem_stage_inst_dmem_ram_69__11_), .D(
        mem_stage_inst_dmem_ram_71__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5304) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1100 ( .A(
        mem_stage_inst_dmem_ram_76__11_), .B(mem_stage_inst_dmem_ram_78__11_), 
        .C(mem_stage_inst_dmem_ram_77__11_), .D(
        mem_stage_inst_dmem_ram_79__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5305) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1099 ( .A(mem_stage_inst_dmem_n5302), 
        .B(mem_stage_inst_dmem_n5303), .C(mem_stage_inst_dmem_n5304), .D(
        mem_stage_inst_dmem_n5305), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5301) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1098 ( .A(
        mem_stage_inst_dmem_ram_192__10_), .B(mem_stage_inst_dmem_ram_194__10_), .C(mem_stage_inst_dmem_ram_193__10_), .D(mem_stage_inst_dmem_ram_195__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5178) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1097 ( .A(
        mem_stage_inst_dmem_ram_196__10_), .B(mem_stage_inst_dmem_ram_198__10_), .C(mem_stage_inst_dmem_ram_197__10_), .D(mem_stage_inst_dmem_ram_199__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5180) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1096 ( .A(
        mem_stage_inst_dmem_ram_204__10_), .B(mem_stage_inst_dmem_ram_206__10_), .C(mem_stage_inst_dmem_ram_205__10_), .D(mem_stage_inst_dmem_ram_207__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5181) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1095 ( .A(mem_stage_inst_dmem_n5178), 
        .B(mem_stage_inst_dmem_n5179), .C(mem_stage_inst_dmem_n5180), .D(
        mem_stage_inst_dmem_n5181), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5177) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1094 ( .A(
        mem_stage_inst_dmem_ram_64__10_), .B(mem_stage_inst_dmem_ram_66__10_), 
        .C(mem_stage_inst_dmem_ram_65__10_), .D(
        mem_stage_inst_dmem_ram_67__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5218) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1093 ( .A(
        mem_stage_inst_dmem_ram_68__10_), .B(mem_stage_inst_dmem_ram_70__10_), 
        .C(mem_stage_inst_dmem_ram_69__10_), .D(
        mem_stage_inst_dmem_ram_71__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5220) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1092 ( .A(
        mem_stage_inst_dmem_ram_76__10_), .B(mem_stage_inst_dmem_ram_78__10_), 
        .C(mem_stage_inst_dmem_ram_77__10_), .D(
        mem_stage_inst_dmem_ram_79__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5221) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1091 ( .A(mem_stage_inst_dmem_n5218), 
        .B(mem_stage_inst_dmem_n5219), .C(mem_stage_inst_dmem_n5220), .D(
        mem_stage_inst_dmem_n5221), .S0(mem_stage_inst_dmem_n215), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5217) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1090 ( .A(
        mem_stage_inst_dmem_ram_192__9_), .B(mem_stage_inst_dmem_ram_194__9_), 
        .C(mem_stage_inst_dmem_ram_193__9_), .D(
        mem_stage_inst_dmem_ram_195__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5094) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1089 ( .A(
        mem_stage_inst_dmem_ram_196__9_), .B(mem_stage_inst_dmem_ram_198__9_), 
        .C(mem_stage_inst_dmem_ram_197__9_), .D(
        mem_stage_inst_dmem_ram_199__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5096) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1088 ( .A(
        mem_stage_inst_dmem_ram_204__9_), .B(mem_stage_inst_dmem_ram_206__9_), 
        .C(mem_stage_inst_dmem_ram_205__9_), .D(
        mem_stage_inst_dmem_ram_207__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5097) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1087 ( .A(mem_stage_inst_dmem_n5094), 
        .B(mem_stage_inst_dmem_n5095), .C(mem_stage_inst_dmem_n5096), .D(
        mem_stage_inst_dmem_n5097), .S0(mem_stage_inst_dmem_n214), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5093) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1086 ( .A(
        mem_stage_inst_dmem_ram_64__9_), .B(mem_stage_inst_dmem_ram_66__9_), 
        .C(mem_stage_inst_dmem_ram_65__9_), .D(mem_stage_inst_dmem_ram_67__9_), 
        .S0(mem_stage_inst_dmem_n147), .S1(ex_pipeline_reg_out[22]), .Y(
        mem_stage_inst_dmem_n5134) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1085 ( .A(
        mem_stage_inst_dmem_ram_68__9_), .B(mem_stage_inst_dmem_ram_70__9_), 
        .C(mem_stage_inst_dmem_ram_69__9_), .D(mem_stage_inst_dmem_ram_71__9_), 
        .S0(mem_stage_inst_dmem_n146), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n5136) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1084 ( .A(
        mem_stage_inst_dmem_ram_76__9_), .B(mem_stage_inst_dmem_ram_78__9_), 
        .C(mem_stage_inst_dmem_ram_77__9_), .D(mem_stage_inst_dmem_ram_79__9_), 
        .S0(mem_stage_inst_dmem_n145), .S1(mem_stage_inst_dmem_n31), .Y(
        mem_stage_inst_dmem_n5137) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1083 ( .A(mem_stage_inst_dmem_n5134), 
        .B(mem_stage_inst_dmem_n5135), .C(mem_stage_inst_dmem_n5136), .D(
        mem_stage_inst_dmem_n5137), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5133) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1082 ( .A(
        mem_stage_inst_dmem_ram_192__8_), .B(mem_stage_inst_dmem_ram_194__8_), 
        .C(mem_stage_inst_dmem_ram_193__8_), .D(
        mem_stage_inst_dmem_ram_195__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5010) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1081 ( .A(
        mem_stage_inst_dmem_ram_196__8_), .B(mem_stage_inst_dmem_ram_198__8_), 
        .C(mem_stage_inst_dmem_ram_197__8_), .D(
        mem_stage_inst_dmem_ram_199__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5012) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1080 ( .A(
        mem_stage_inst_dmem_ram_204__8_), .B(mem_stage_inst_dmem_ram_206__8_), 
        .C(mem_stage_inst_dmem_ram_205__8_), .D(
        mem_stage_inst_dmem_ram_207__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5013) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1079 ( .A(mem_stage_inst_dmem_n5010), 
        .B(mem_stage_inst_dmem_n5011), .C(mem_stage_inst_dmem_n5012), .D(
        mem_stage_inst_dmem_n5013), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5009) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1078 ( .A(
        mem_stage_inst_dmem_ram_64__8_), .B(mem_stage_inst_dmem_ram_66__8_), 
        .C(mem_stage_inst_dmem_ram_65__8_), .D(mem_stage_inst_dmem_ram_67__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5050) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1077 ( .A(
        mem_stage_inst_dmem_ram_68__8_), .B(mem_stage_inst_dmem_ram_70__8_), 
        .C(mem_stage_inst_dmem_ram_69__8_), .D(mem_stage_inst_dmem_ram_71__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5052) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1076 ( .A(
        mem_stage_inst_dmem_ram_76__8_), .B(mem_stage_inst_dmem_ram_78__8_), 
        .C(mem_stage_inst_dmem_ram_77__8_), .D(mem_stage_inst_dmem_ram_79__8_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n14), .Y(
        mem_stage_inst_dmem_n5053) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1075 ( .A(mem_stage_inst_dmem_n5050), 
        .B(mem_stage_inst_dmem_n5051), .C(mem_stage_inst_dmem_n5052), .D(
        mem_stage_inst_dmem_n5053), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5049) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1074 ( .A(
        mem_stage_inst_dmem_ram_192__7_), .B(mem_stage_inst_dmem_ram_194__7_), 
        .C(mem_stage_inst_dmem_ram_193__7_), .D(
        mem_stage_inst_dmem_ram_195__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4926) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1073 ( .A(
        mem_stage_inst_dmem_ram_196__7_), .B(mem_stage_inst_dmem_ram_198__7_), 
        .C(mem_stage_inst_dmem_ram_197__7_), .D(
        mem_stage_inst_dmem_ram_199__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4928) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1072 ( .A(
        mem_stage_inst_dmem_ram_204__7_), .B(mem_stage_inst_dmem_ram_206__7_), 
        .C(mem_stage_inst_dmem_ram_205__7_), .D(
        mem_stage_inst_dmem_ram_207__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4929) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1071 ( .A(mem_stage_inst_dmem_n4926), 
        .B(mem_stage_inst_dmem_n4927), .C(mem_stage_inst_dmem_n4928), .D(
        mem_stage_inst_dmem_n4929), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4925) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1070 ( .A(
        mem_stage_inst_dmem_ram_64__7_), .B(mem_stage_inst_dmem_ram_66__7_), 
        .C(mem_stage_inst_dmem_ram_65__7_), .D(mem_stage_inst_dmem_ram_67__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4966) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1069 ( .A(
        mem_stage_inst_dmem_ram_68__7_), .B(mem_stage_inst_dmem_ram_70__7_), 
        .C(mem_stage_inst_dmem_ram_69__7_), .D(mem_stage_inst_dmem_ram_71__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4968) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1068 ( .A(
        mem_stage_inst_dmem_ram_76__7_), .B(mem_stage_inst_dmem_ram_78__7_), 
        .C(mem_stage_inst_dmem_ram_77__7_), .D(mem_stage_inst_dmem_ram_79__7_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n4969) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1067 ( .A(mem_stage_inst_dmem_n4966), 
        .B(mem_stage_inst_dmem_n4967), .C(mem_stage_inst_dmem_n4968), .D(
        mem_stage_inst_dmem_n4969), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4965) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1066 ( .A(
        mem_stage_inst_dmem_ram_192__6_), .B(mem_stage_inst_dmem_ram_194__6_), 
        .C(mem_stage_inst_dmem_ram_193__6_), .D(
        mem_stage_inst_dmem_ram_195__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4842) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1065 ( .A(
        mem_stage_inst_dmem_ram_196__6_), .B(mem_stage_inst_dmem_ram_198__6_), 
        .C(mem_stage_inst_dmem_ram_197__6_), .D(
        mem_stage_inst_dmem_ram_199__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4844) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1064 ( .A(
        mem_stage_inst_dmem_ram_204__6_), .B(mem_stage_inst_dmem_ram_206__6_), 
        .C(mem_stage_inst_dmem_ram_205__6_), .D(
        mem_stage_inst_dmem_ram_207__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4845) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1063 ( .A(mem_stage_inst_dmem_n4842), 
        .B(mem_stage_inst_dmem_n4843), .C(mem_stage_inst_dmem_n4844), .D(
        mem_stage_inst_dmem_n4845), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4841) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1062 ( .A(
        mem_stage_inst_dmem_ram_64__6_), .B(mem_stage_inst_dmem_ram_66__6_), 
        .C(mem_stage_inst_dmem_ram_65__6_), .D(mem_stage_inst_dmem_ram_67__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4882) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1061 ( .A(
        mem_stage_inst_dmem_ram_68__6_), .B(mem_stage_inst_dmem_ram_70__6_), 
        .C(mem_stage_inst_dmem_ram_69__6_), .D(mem_stage_inst_dmem_ram_71__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4884) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1060 ( .A(
        mem_stage_inst_dmem_ram_76__6_), .B(mem_stage_inst_dmem_ram_78__6_), 
        .C(mem_stage_inst_dmem_ram_77__6_), .D(mem_stage_inst_dmem_ram_79__6_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n4885) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1059 ( .A(mem_stage_inst_dmem_n4882), 
        .B(mem_stage_inst_dmem_n4883), .C(mem_stage_inst_dmem_n4884), .D(
        mem_stage_inst_dmem_n4885), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4881) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1058 ( .A(
        mem_stage_inst_dmem_ram_192__5_), .B(mem_stage_inst_dmem_ram_194__5_), 
        .C(mem_stage_inst_dmem_ram_193__5_), .D(
        mem_stage_inst_dmem_ram_195__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4758) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1057 ( .A(
        mem_stage_inst_dmem_ram_196__5_), .B(mem_stage_inst_dmem_ram_198__5_), 
        .C(mem_stage_inst_dmem_ram_197__5_), .D(
        mem_stage_inst_dmem_ram_199__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4760) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1056 ( .A(
        mem_stage_inst_dmem_ram_204__5_), .B(mem_stage_inst_dmem_ram_206__5_), 
        .C(mem_stage_inst_dmem_ram_205__5_), .D(
        mem_stage_inst_dmem_ram_207__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4761) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1055 ( .A(mem_stage_inst_dmem_n4758), 
        .B(mem_stage_inst_dmem_n4759), .C(mem_stage_inst_dmem_n4760), .D(
        mem_stage_inst_dmem_n4761), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4757) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1054 ( .A(
        mem_stage_inst_dmem_ram_64__5_), .B(mem_stage_inst_dmem_ram_66__5_), 
        .C(mem_stage_inst_dmem_ram_65__5_), .D(mem_stage_inst_dmem_ram_67__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4798) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1053 ( .A(
        mem_stage_inst_dmem_ram_68__5_), .B(mem_stage_inst_dmem_ram_70__5_), 
        .C(mem_stage_inst_dmem_ram_69__5_), .D(mem_stage_inst_dmem_ram_71__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4800) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1052 ( .A(
        mem_stage_inst_dmem_ram_76__5_), .B(mem_stage_inst_dmem_ram_78__5_), 
        .C(mem_stage_inst_dmem_ram_77__5_), .D(mem_stage_inst_dmem_ram_79__5_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n4801) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1051 ( .A(mem_stage_inst_dmem_n4798), 
        .B(mem_stage_inst_dmem_n4799), .C(mem_stage_inst_dmem_n4800), .D(
        mem_stage_inst_dmem_n4801), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4797) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1050 ( .A(
        mem_stage_inst_dmem_ram_192__4_), .B(mem_stage_inst_dmem_ram_194__4_), 
        .C(mem_stage_inst_dmem_ram_193__4_), .D(
        mem_stage_inst_dmem_ram_195__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4674) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1049 ( .A(
        mem_stage_inst_dmem_ram_196__4_), .B(mem_stage_inst_dmem_ram_198__4_), 
        .C(mem_stage_inst_dmem_ram_197__4_), .D(
        mem_stage_inst_dmem_ram_199__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4676) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1048 ( .A(
        mem_stage_inst_dmem_ram_204__4_), .B(mem_stage_inst_dmem_ram_206__4_), 
        .C(mem_stage_inst_dmem_ram_205__4_), .D(
        mem_stage_inst_dmem_ram_207__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4677) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1047 ( .A(mem_stage_inst_dmem_n4674), 
        .B(mem_stage_inst_dmem_n4675), .C(mem_stage_inst_dmem_n4676), .D(
        mem_stage_inst_dmem_n4677), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4673) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1046 ( .A(
        mem_stage_inst_dmem_ram_64__4_), .B(mem_stage_inst_dmem_ram_66__4_), 
        .C(mem_stage_inst_dmem_ram_65__4_), .D(mem_stage_inst_dmem_ram_67__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4714) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1045 ( .A(
        mem_stage_inst_dmem_ram_68__4_), .B(mem_stage_inst_dmem_ram_70__4_), 
        .C(mem_stage_inst_dmem_ram_69__4_), .D(mem_stage_inst_dmem_ram_71__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4716) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1044 ( .A(
        mem_stage_inst_dmem_ram_76__4_), .B(mem_stage_inst_dmem_ram_78__4_), 
        .C(mem_stage_inst_dmem_ram_77__4_), .D(mem_stage_inst_dmem_ram_79__4_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n4717) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1043 ( .A(mem_stage_inst_dmem_n4714), 
        .B(mem_stage_inst_dmem_n4715), .C(mem_stage_inst_dmem_n4716), .D(
        mem_stage_inst_dmem_n4717), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4713) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1042 ( .A(
        mem_stage_inst_dmem_ram_192__3_), .B(mem_stage_inst_dmem_ram_194__3_), 
        .C(mem_stage_inst_dmem_ram_193__3_), .D(
        mem_stage_inst_dmem_ram_195__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n494) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1041 ( .A(
        mem_stage_inst_dmem_ram_196__3_), .B(mem_stage_inst_dmem_ram_198__3_), 
        .C(mem_stage_inst_dmem_ram_197__3_), .D(
        mem_stage_inst_dmem_ram_199__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n496) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1040 ( .A(
        mem_stage_inst_dmem_ram_204__3_), .B(mem_stage_inst_dmem_ram_206__3_), 
        .C(mem_stage_inst_dmem_ram_205__3_), .D(
        mem_stage_inst_dmem_ram_207__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n497) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1039 ( .A(mem_stage_inst_dmem_n494), 
        .B(mem_stage_inst_dmem_n495), .C(mem_stage_inst_dmem_n496), .D(
        mem_stage_inst_dmem_n497), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n493) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1038 ( .A(
        mem_stage_inst_dmem_ram_64__3_), .B(mem_stage_inst_dmem_ram_66__3_), 
        .C(mem_stage_inst_dmem_ram_65__3_), .D(mem_stage_inst_dmem_ram_67__3_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n534) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1037 ( .A(
        mem_stage_inst_dmem_ram_68__3_), .B(mem_stage_inst_dmem_ram_70__3_), 
        .C(mem_stage_inst_dmem_ram_69__3_), .D(mem_stage_inst_dmem_ram_71__3_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n536) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1036 ( .A(
        mem_stage_inst_dmem_ram_76__3_), .B(mem_stage_inst_dmem_ram_78__3_), 
        .C(mem_stage_inst_dmem_ram_77__3_), .D(mem_stage_inst_dmem_ram_79__3_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n537) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1035 ( .A(mem_stage_inst_dmem_n534), 
        .B(mem_stage_inst_dmem_n535), .C(mem_stage_inst_dmem_n536), .D(
        mem_stage_inst_dmem_n537), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n533) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1034 ( .A(
        mem_stage_inst_dmem_ram_192__2_), .B(mem_stage_inst_dmem_ram_194__2_), 
        .C(mem_stage_inst_dmem_ram_193__2_), .D(
        mem_stage_inst_dmem_ram_195__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n410) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1033 ( .A(
        mem_stage_inst_dmem_ram_196__2_), .B(mem_stage_inst_dmem_ram_198__2_), 
        .C(mem_stage_inst_dmem_ram_197__2_), .D(
        mem_stage_inst_dmem_ram_199__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n412) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1032 ( .A(
        mem_stage_inst_dmem_ram_204__2_), .B(mem_stage_inst_dmem_ram_206__2_), 
        .C(mem_stage_inst_dmem_ram_205__2_), .D(
        mem_stage_inst_dmem_ram_207__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n413) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1031 ( .A(mem_stage_inst_dmem_n410), 
        .B(mem_stage_inst_dmem_n411), .C(mem_stage_inst_dmem_n412), .D(
        mem_stage_inst_dmem_n413), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n409) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1030 ( .A(
        mem_stage_inst_dmem_ram_64__2_), .B(mem_stage_inst_dmem_ram_66__2_), 
        .C(mem_stage_inst_dmem_ram_65__2_), .D(mem_stage_inst_dmem_ram_67__2_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n450) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1029 ( .A(
        mem_stage_inst_dmem_ram_68__2_), .B(mem_stage_inst_dmem_ram_70__2_), 
        .C(mem_stage_inst_dmem_ram_69__2_), .D(mem_stage_inst_dmem_ram_71__2_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n452) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1028 ( .A(
        mem_stage_inst_dmem_ram_76__2_), .B(mem_stage_inst_dmem_ram_78__2_), 
        .C(mem_stage_inst_dmem_ram_77__2_), .D(mem_stage_inst_dmem_ram_79__2_), 
        .S0(mem_stage_inst_dmem_n128), .S1(mem_stage_inst_dmem_n30), .Y(
        mem_stage_inst_dmem_n453) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1027 ( .A(mem_stage_inst_dmem_n450), 
        .B(mem_stage_inst_dmem_n451), .C(mem_stage_inst_dmem_n452), .D(
        mem_stage_inst_dmem_n453), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n449) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1026 ( .A(
        mem_stage_inst_dmem_ram_192__1_), .B(mem_stage_inst_dmem_ram_194__1_), 
        .C(mem_stage_inst_dmem_ram_193__1_), .D(
        mem_stage_inst_dmem_ram_195__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n326) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1025 ( .A(
        mem_stage_inst_dmem_ram_196__1_), .B(mem_stage_inst_dmem_ram_198__1_), 
        .C(mem_stage_inst_dmem_ram_197__1_), .D(
        mem_stage_inst_dmem_ram_199__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n328) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1024 ( .A(
        mem_stage_inst_dmem_ram_204__1_), .B(mem_stage_inst_dmem_ram_206__1_), 
        .C(mem_stage_inst_dmem_ram_205__1_), .D(
        mem_stage_inst_dmem_ram_207__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n329) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1023 ( .A(mem_stage_inst_dmem_n326), 
        .B(mem_stage_inst_dmem_n327), .C(mem_stage_inst_dmem_n328), .D(
        mem_stage_inst_dmem_n329), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n325) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1022 ( .A(
        mem_stage_inst_dmem_ram_64__1_), .B(mem_stage_inst_dmem_ram_66__1_), 
        .C(mem_stage_inst_dmem_ram_65__1_), .D(mem_stage_inst_dmem_ram_67__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n366) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1021 ( .A(
        mem_stage_inst_dmem_ram_68__1_), .B(mem_stage_inst_dmem_ram_70__1_), 
        .C(mem_stage_inst_dmem_ram_69__1_), .D(mem_stage_inst_dmem_ram_71__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n368) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1020 ( .A(
        mem_stage_inst_dmem_ram_76__1_), .B(mem_stage_inst_dmem_ram_78__1_), 
        .C(mem_stage_inst_dmem_ram_77__1_), .D(mem_stage_inst_dmem_ram_79__1_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n45), .Y(
        mem_stage_inst_dmem_n369) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1019 ( .A(mem_stage_inst_dmem_n366), 
        .B(mem_stage_inst_dmem_n367), .C(mem_stage_inst_dmem_n368), .D(
        mem_stage_inst_dmem_n369), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n365) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1018 ( .A(
        mem_stage_inst_dmem_ram_192__0_), .B(mem_stage_inst_dmem_ram_194__0_), 
        .C(mem_stage_inst_dmem_ram_193__0_), .D(
        mem_stage_inst_dmem_ram_195__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n242) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1017 ( .A(
        mem_stage_inst_dmem_ram_196__0_), .B(mem_stage_inst_dmem_ram_198__0_), 
        .C(mem_stage_inst_dmem_ram_197__0_), .D(
        mem_stage_inst_dmem_ram_199__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n244) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1016 ( .A(
        mem_stage_inst_dmem_ram_204__0_), .B(mem_stage_inst_dmem_ram_206__0_), 
        .C(mem_stage_inst_dmem_ram_205__0_), .D(
        mem_stage_inst_dmem_ram_207__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n245) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1015 ( .A(mem_stage_inst_dmem_n242), 
        .B(mem_stage_inst_dmem_n243), .C(mem_stage_inst_dmem_n244), .D(
        mem_stage_inst_dmem_n245), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n241) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1014 ( .A(
        mem_stage_inst_dmem_ram_64__0_), .B(mem_stage_inst_dmem_ram_66__0_), 
        .C(mem_stage_inst_dmem_ram_65__0_), .D(mem_stage_inst_dmem_ram_67__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n282) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1013 ( .A(
        mem_stage_inst_dmem_ram_68__0_), .B(mem_stage_inst_dmem_ram_70__0_), 
        .C(mem_stage_inst_dmem_ram_69__0_), .D(mem_stage_inst_dmem_ram_71__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n284) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1012 ( .A(
        mem_stage_inst_dmem_ram_76__0_), .B(mem_stage_inst_dmem_ram_78__0_), 
        .C(mem_stage_inst_dmem_ram_77__0_), .D(mem_stage_inst_dmem_ram_79__0_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n40), .Y(
        mem_stage_inst_dmem_n285) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1011 ( .A(mem_stage_inst_dmem_n282), 
        .B(mem_stage_inst_dmem_n283), .C(mem_stage_inst_dmem_n284), .D(
        mem_stage_inst_dmem_n285), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n281) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1010 ( .A(
        mem_stage_inst_dmem_ram_48__15_), .B(mem_stage_inst_dmem_ram_50__15_), 
        .C(mem_stage_inst_dmem_ram_49__15_), .D(
        mem_stage_inst_dmem_ram_51__15_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n5643) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1009 ( .A(
        mem_stage_inst_dmem_ram_16__15_), .B(mem_stage_inst_dmem_ram_18__15_), 
        .C(mem_stage_inst_dmem_ram_17__15_), .D(
        mem_stage_inst_dmem_ram_19__15_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n5653) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1008 ( .A(
        mem_stage_inst_dmem_ram_0__15_), .B(mem_stage_inst_dmem_ram_2__15_), 
        .C(mem_stage_inst_dmem_ram_1__15_), .D(mem_stage_inst_dmem_ram_3__15_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n65), .Y(
        mem_stage_inst_dmem_n5658) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1007 ( .A(
        mem_stage_inst_dmem_ram_176__15_), .B(mem_stage_inst_dmem_ram_178__15_), .C(mem_stage_inst_dmem_ram_177__15_), .D(mem_stage_inst_dmem_ram_179__15_), 
        .S0(mem_stage_inst_dmem_n155), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5603) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1006 ( .A(
        mem_stage_inst_dmem_ram_144__15_), .B(mem_stage_inst_dmem_ram_146__15_), .C(mem_stage_inst_dmem_ram_145__15_), .D(mem_stage_inst_dmem_ram_147__15_), 
        .S0(mem_stage_inst_dmem_n156), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5613) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1005 ( .A(
        mem_stage_inst_dmem_ram_128__15_), .B(mem_stage_inst_dmem_ram_130__15_), .C(mem_stage_inst_dmem_ram_129__15_), .D(mem_stage_inst_dmem_ram_131__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n37), .Y(
        mem_stage_inst_dmem_n5618) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1004 ( .A(
        mem_stage_inst_dmem_ram_48__14_), .B(mem_stage_inst_dmem_ram_50__14_), 
        .C(mem_stage_inst_dmem_ram_49__14_), .D(
        mem_stage_inst_dmem_ram_51__14_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5559) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1003 ( .A(
        mem_stage_inst_dmem_ram_16__14_), .B(mem_stage_inst_dmem_ram_18__14_), 
        .C(mem_stage_inst_dmem_ram_17__14_), .D(
        mem_stage_inst_dmem_ram_19__14_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5569) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1002 ( .A(
        mem_stage_inst_dmem_ram_0__14_), .B(mem_stage_inst_dmem_ram_2__14_), 
        .C(mem_stage_inst_dmem_ram_1__14_), .D(mem_stage_inst_dmem_ram_3__14_), 
        .S0(mem_stage_inst_dmem_n141), .S1(mem_stage_inst_dmem_n28), .Y(
        mem_stage_inst_dmem_n5574) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1001 ( .A(
        mem_stage_inst_dmem_ram_176__14_), .B(mem_stage_inst_dmem_ram_178__14_), .C(mem_stage_inst_dmem_ram_177__14_), .D(mem_stage_inst_dmem_ram_179__14_), 
        .S0(mem_stage_inst_dmem_n111), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5519) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u1000 ( .A(
        mem_stage_inst_dmem_ram_144__14_), .B(mem_stage_inst_dmem_ram_146__14_), .C(mem_stage_inst_dmem_ram_145__14_), .D(mem_stage_inst_dmem_ram_147__14_), 
        .S0(mem_stage_inst_dmem_n112), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5529) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u999 ( .A(
        mem_stage_inst_dmem_ram_128__14_), .B(mem_stage_inst_dmem_ram_130__14_), .C(mem_stage_inst_dmem_ram_129__14_), .D(mem_stage_inst_dmem_ram_131__14_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5534) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u998 ( .A(
        mem_stage_inst_dmem_ram_48__13_), .B(mem_stage_inst_dmem_ram_50__13_), 
        .C(mem_stage_inst_dmem_ram_49__13_), .D(
        mem_stage_inst_dmem_ram_51__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5475) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u997 ( .A(
        mem_stage_inst_dmem_ram_16__13_), .B(mem_stage_inst_dmem_ram_18__13_), 
        .C(mem_stage_inst_dmem_ram_17__13_), .D(
        mem_stage_inst_dmem_ram_19__13_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n5485) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u996 ( .A(mem_stage_inst_dmem_ram_0__13_), .B(mem_stage_inst_dmem_ram_2__13_), .C(mem_stage_inst_dmem_ram_1__13_), .D(
        mem_stage_inst_dmem_ram_3__13_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n5490) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u995 ( .A(
        mem_stage_inst_dmem_ram_176__13_), .B(mem_stage_inst_dmem_ram_178__13_), .C(mem_stage_inst_dmem_ram_177__13_), .D(mem_stage_inst_dmem_ram_179__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(ex_pipeline_reg_out[22]), .Y(
        mem_stage_inst_dmem_n5435) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u994 ( .A(
        mem_stage_inst_dmem_ram_144__13_), .B(mem_stage_inst_dmem_ram_146__13_), .C(mem_stage_inst_dmem_ram_145__13_), .D(mem_stage_inst_dmem_ram_147__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5445) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u993 ( .A(
        mem_stage_inst_dmem_ram_128__13_), .B(mem_stage_inst_dmem_ram_130__13_), .C(mem_stage_inst_dmem_ram_129__13_), .D(mem_stage_inst_dmem_ram_131__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5450) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u992 ( .A(
        mem_stage_inst_dmem_ram_48__12_), .B(mem_stage_inst_dmem_ram_50__12_), 
        .C(mem_stage_inst_dmem_ram_49__12_), .D(
        mem_stage_inst_dmem_ram_51__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n5391) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u991 ( .A(
        mem_stage_inst_dmem_ram_16__12_), .B(mem_stage_inst_dmem_ram_18__12_), 
        .C(mem_stage_inst_dmem_ram_17__12_), .D(
        mem_stage_inst_dmem_ram_19__12_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5401) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u990 ( .A(mem_stage_inst_dmem_ram_0__12_), .B(mem_stage_inst_dmem_ram_2__12_), .C(mem_stage_inst_dmem_ram_1__12_), .D(
        mem_stage_inst_dmem_ram_3__12_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5406) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u989 ( .A(
        mem_stage_inst_dmem_ram_176__12_), .B(mem_stage_inst_dmem_ram_178__12_), .C(mem_stage_inst_dmem_ram_177__12_), .D(mem_stage_inst_dmem_ram_179__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5351) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u988 ( .A(
        mem_stage_inst_dmem_ram_144__12_), .B(mem_stage_inst_dmem_ram_146__12_), .C(mem_stage_inst_dmem_ram_145__12_), .D(mem_stage_inst_dmem_ram_147__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5361) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u987 ( .A(
        mem_stage_inst_dmem_ram_128__12_), .B(mem_stage_inst_dmem_ram_130__12_), .C(mem_stage_inst_dmem_ram_129__12_), .D(mem_stage_inst_dmem_ram_131__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5366) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u986 ( .A(
        mem_stage_inst_dmem_ram_48__11_), .B(mem_stage_inst_dmem_ram_50__11_), 
        .C(mem_stage_inst_dmem_ram_49__11_), .D(
        mem_stage_inst_dmem_ram_51__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5307) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u985 ( .A(
        mem_stage_inst_dmem_ram_16__11_), .B(mem_stage_inst_dmem_ram_18__11_), 
        .C(mem_stage_inst_dmem_ram_17__11_), .D(
        mem_stage_inst_dmem_ram_19__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5317) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u984 ( .A(mem_stage_inst_dmem_ram_0__11_), .B(mem_stage_inst_dmem_ram_2__11_), .C(mem_stage_inst_dmem_ram_1__11_), .D(
        mem_stage_inst_dmem_ram_3__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5322) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u983 ( .A(
        mem_stage_inst_dmem_ram_176__11_), .B(mem_stage_inst_dmem_ram_178__11_), .C(mem_stage_inst_dmem_ram_177__11_), .D(mem_stage_inst_dmem_ram_179__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5267) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u982 ( .A(
        mem_stage_inst_dmem_ram_144__11_), .B(mem_stage_inst_dmem_ram_146__11_), .C(mem_stage_inst_dmem_ram_145__11_), .D(mem_stage_inst_dmem_ram_147__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5277) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u981 ( .A(
        mem_stage_inst_dmem_ram_128__11_), .B(mem_stage_inst_dmem_ram_130__11_), .C(mem_stage_inst_dmem_ram_129__11_), .D(mem_stage_inst_dmem_ram_131__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5282) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u980 ( .A(
        mem_stage_inst_dmem_ram_48__10_), .B(mem_stage_inst_dmem_ram_50__10_), 
        .C(mem_stage_inst_dmem_ram_49__10_), .D(
        mem_stage_inst_dmem_ram_51__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5223) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u979 ( .A(
        mem_stage_inst_dmem_ram_16__10_), .B(mem_stage_inst_dmem_ram_18__10_), 
        .C(mem_stage_inst_dmem_ram_17__10_), .D(
        mem_stage_inst_dmem_ram_19__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5233) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u978 ( .A(mem_stage_inst_dmem_ram_0__10_), .B(mem_stage_inst_dmem_ram_2__10_), .C(mem_stage_inst_dmem_ram_1__10_), .D(
        mem_stage_inst_dmem_ram_3__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5238) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u977 ( .A(
        mem_stage_inst_dmem_ram_176__10_), .B(mem_stage_inst_dmem_ram_178__10_), .C(mem_stage_inst_dmem_ram_177__10_), .D(mem_stage_inst_dmem_ram_179__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5183) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u976 ( .A(
        mem_stage_inst_dmem_ram_144__10_), .B(mem_stage_inst_dmem_ram_146__10_), .C(mem_stage_inst_dmem_ram_145__10_), .D(mem_stage_inst_dmem_ram_147__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5193) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u975 ( .A(
        mem_stage_inst_dmem_ram_128__10_), .B(mem_stage_inst_dmem_ram_130__10_), .C(mem_stage_inst_dmem_ram_129__10_), .D(mem_stage_inst_dmem_ram_131__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5198) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u974 ( .A(mem_stage_inst_dmem_ram_48__9_), .B(mem_stage_inst_dmem_ram_50__9_), .C(mem_stage_inst_dmem_ram_49__9_), .D(
        mem_stage_inst_dmem_ram_51__9_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5139) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u973 ( .A(mem_stage_inst_dmem_ram_16__9_), .B(mem_stage_inst_dmem_ram_18__9_), .C(mem_stage_inst_dmem_ram_17__9_), .D(
        mem_stage_inst_dmem_ram_19__9_), .S0(mem_stage_inst_dmem_n101), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n5149) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u972 ( .A(mem_stage_inst_dmem_ram_0__9_), 
        .B(mem_stage_inst_dmem_ram_2__9_), .C(mem_stage_inst_dmem_ram_1__9_), 
        .D(mem_stage_inst_dmem_ram_3__9_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n5154) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u971 ( .A(
        mem_stage_inst_dmem_ram_176__9_), .B(mem_stage_inst_dmem_ram_178__9_), 
        .C(mem_stage_inst_dmem_ram_177__9_), .D(
        mem_stage_inst_dmem_ram_179__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5099) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u970 ( .A(
        mem_stage_inst_dmem_ram_144__9_), .B(mem_stage_inst_dmem_ram_146__9_), 
        .C(mem_stage_inst_dmem_ram_145__9_), .D(
        mem_stage_inst_dmem_ram_147__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5109) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u969 ( .A(
        mem_stage_inst_dmem_ram_128__9_), .B(mem_stage_inst_dmem_ram_130__9_), 
        .C(mem_stage_inst_dmem_ram_129__9_), .D(
        mem_stage_inst_dmem_ram_131__9_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5114) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u968 ( .A(mem_stage_inst_dmem_ram_48__8_), .B(mem_stage_inst_dmem_ram_50__8_), .C(mem_stage_inst_dmem_ram_49__8_), .D(
        mem_stage_inst_dmem_ram_51__8_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5055) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u967 ( .A(mem_stage_inst_dmem_ram_16__8_), .B(mem_stage_inst_dmem_ram_18__8_), .C(mem_stage_inst_dmem_ram_17__8_), .D(
        mem_stage_inst_dmem_ram_19__8_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5065) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u966 ( .A(mem_stage_inst_dmem_ram_0__8_), 
        .B(mem_stage_inst_dmem_ram_2__8_), .C(mem_stage_inst_dmem_ram_1__8_), 
        .D(mem_stage_inst_dmem_ram_3__8_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5070) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u965 ( .A(
        mem_stage_inst_dmem_ram_176__8_), .B(mem_stage_inst_dmem_ram_178__8_), 
        .C(mem_stage_inst_dmem_ram_177__8_), .D(
        mem_stage_inst_dmem_ram_179__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5015) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u964 ( .A(
        mem_stage_inst_dmem_ram_144__8_), .B(mem_stage_inst_dmem_ram_146__8_), 
        .C(mem_stage_inst_dmem_ram_145__8_), .D(
        mem_stage_inst_dmem_ram_147__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5025) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u963 ( .A(
        mem_stage_inst_dmem_ram_128__8_), .B(mem_stage_inst_dmem_ram_130__8_), 
        .C(mem_stage_inst_dmem_ram_129__8_), .D(
        mem_stage_inst_dmem_ram_131__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5030) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u962 ( .A(mem_stage_inst_dmem_ram_48__7_), .B(mem_stage_inst_dmem_ram_50__7_), .C(mem_stage_inst_dmem_ram_49__7_), .D(
        mem_stage_inst_dmem_ram_51__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4971) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u961 ( .A(mem_stage_inst_dmem_ram_16__7_), .B(mem_stage_inst_dmem_ram_18__7_), .C(mem_stage_inst_dmem_ram_17__7_), .D(
        mem_stage_inst_dmem_ram_19__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4981) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u960 ( .A(mem_stage_inst_dmem_ram_0__7_), 
        .B(mem_stage_inst_dmem_ram_2__7_), .C(mem_stage_inst_dmem_ram_1__7_), 
        .D(mem_stage_inst_dmem_ram_3__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4986) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u959 ( .A(
        mem_stage_inst_dmem_ram_176__7_), .B(mem_stage_inst_dmem_ram_178__7_), 
        .C(mem_stage_inst_dmem_ram_177__7_), .D(
        mem_stage_inst_dmem_ram_179__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4931) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u958 ( .A(
        mem_stage_inst_dmem_ram_144__7_), .B(mem_stage_inst_dmem_ram_146__7_), 
        .C(mem_stage_inst_dmem_ram_145__7_), .D(
        mem_stage_inst_dmem_ram_147__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4941) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u957 ( .A(
        mem_stage_inst_dmem_ram_128__7_), .B(mem_stage_inst_dmem_ram_130__7_), 
        .C(mem_stage_inst_dmem_ram_129__7_), .D(
        mem_stage_inst_dmem_ram_131__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4946) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u956 ( .A(mem_stage_inst_dmem_ram_48__6_), .B(mem_stage_inst_dmem_ram_50__6_), .C(mem_stage_inst_dmem_ram_49__6_), .D(
        mem_stage_inst_dmem_ram_51__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4887) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u955 ( .A(mem_stage_inst_dmem_ram_16__6_), .B(mem_stage_inst_dmem_ram_18__6_), .C(mem_stage_inst_dmem_ram_17__6_), .D(
        mem_stage_inst_dmem_ram_19__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4897) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u954 ( .A(mem_stage_inst_dmem_ram_0__6_), 
        .B(mem_stage_inst_dmem_ram_2__6_), .C(mem_stage_inst_dmem_ram_1__6_), 
        .D(mem_stage_inst_dmem_ram_3__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4902) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u953 ( .A(
        mem_stage_inst_dmem_ram_176__6_), .B(mem_stage_inst_dmem_ram_178__6_), 
        .C(mem_stage_inst_dmem_ram_177__6_), .D(
        mem_stage_inst_dmem_ram_179__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4847) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u952 ( .A(
        mem_stage_inst_dmem_ram_144__6_), .B(mem_stage_inst_dmem_ram_146__6_), 
        .C(mem_stage_inst_dmem_ram_145__6_), .D(
        mem_stage_inst_dmem_ram_147__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4857) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u951 ( .A(
        mem_stage_inst_dmem_ram_128__6_), .B(mem_stage_inst_dmem_ram_130__6_), 
        .C(mem_stage_inst_dmem_ram_129__6_), .D(
        mem_stage_inst_dmem_ram_131__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4862) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u950 ( .A(mem_stage_inst_dmem_ram_48__5_), .B(mem_stage_inst_dmem_ram_50__5_), .C(mem_stage_inst_dmem_ram_49__5_), .D(
        mem_stage_inst_dmem_ram_51__5_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n4803) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u949 ( .A(mem_stage_inst_dmem_ram_16__5_), .B(mem_stage_inst_dmem_ram_18__5_), .C(mem_stage_inst_dmem_ram_17__5_), .D(
        mem_stage_inst_dmem_ram_19__5_), .S0(mem_stage_inst_dmem_n164), .S1(
        ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4813) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u948 ( .A(mem_stage_inst_dmem_ram_0__5_), 
        .B(mem_stage_inst_dmem_ram_2__5_), .C(mem_stage_inst_dmem_ram_1__5_), 
        .D(mem_stage_inst_dmem_ram_3__5_), .S0(mem_stage_inst_dmem_n164), .S1(
        ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4818) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u947 ( .A(
        mem_stage_inst_dmem_ram_176__5_), .B(mem_stage_inst_dmem_ram_178__5_), 
        .C(mem_stage_inst_dmem_ram_177__5_), .D(
        mem_stage_inst_dmem_ram_179__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4763) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u946 ( .A(
        mem_stage_inst_dmem_ram_144__5_), .B(mem_stage_inst_dmem_ram_146__5_), 
        .C(mem_stage_inst_dmem_ram_145__5_), .D(
        mem_stage_inst_dmem_ram_147__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4773) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u945 ( .A(
        mem_stage_inst_dmem_ram_128__5_), .B(mem_stage_inst_dmem_ram_130__5_), 
        .C(mem_stage_inst_dmem_ram_129__5_), .D(
        mem_stage_inst_dmem_ram_131__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4778) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u944 ( .A(mem_stage_inst_dmem_ram_48__4_), .B(mem_stage_inst_dmem_ram_50__4_), .C(mem_stage_inst_dmem_ram_49__4_), .D(
        mem_stage_inst_dmem_ram_51__4_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n4719) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u943 ( .A(mem_stage_inst_dmem_ram_16__4_), .B(mem_stage_inst_dmem_ram_18__4_), .C(mem_stage_inst_dmem_ram_17__4_), .D(
        mem_stage_inst_dmem_ram_19__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4729) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u942 ( .A(mem_stage_inst_dmem_ram_0__4_), 
        .B(mem_stage_inst_dmem_ram_2__4_), .C(mem_stage_inst_dmem_ram_1__4_), 
        .D(mem_stage_inst_dmem_ram_3__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4734) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u941 ( .A(
        mem_stage_inst_dmem_ram_176__4_), .B(mem_stage_inst_dmem_ram_178__4_), 
        .C(mem_stage_inst_dmem_ram_177__4_), .D(
        mem_stage_inst_dmem_ram_179__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4679) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u940 ( .A(
        mem_stage_inst_dmem_ram_144__4_), .B(mem_stage_inst_dmem_ram_146__4_), 
        .C(mem_stage_inst_dmem_ram_145__4_), .D(
        mem_stage_inst_dmem_ram_147__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4689) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u939 ( .A(
        mem_stage_inst_dmem_ram_128__4_), .B(mem_stage_inst_dmem_ram_130__4_), 
        .C(mem_stage_inst_dmem_ram_129__4_), .D(
        mem_stage_inst_dmem_ram_131__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4694) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u938 ( .A(mem_stage_inst_dmem_ram_48__3_), .B(mem_stage_inst_dmem_ram_50__3_), .C(mem_stage_inst_dmem_ram_49__3_), .D(
        mem_stage_inst_dmem_ram_51__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n539) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u937 ( .A(mem_stage_inst_dmem_ram_16__3_), .B(mem_stage_inst_dmem_ram_18__3_), .C(mem_stage_inst_dmem_ram_17__3_), .D(
        mem_stage_inst_dmem_ram_19__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n549) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u936 ( .A(mem_stage_inst_dmem_ram_0__3_), 
        .B(mem_stage_inst_dmem_ram_2__3_), .C(mem_stage_inst_dmem_ram_1__3_), 
        .D(mem_stage_inst_dmem_ram_3__3_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n554) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u935 ( .A(
        mem_stage_inst_dmem_ram_176__3_), .B(mem_stage_inst_dmem_ram_178__3_), 
        .C(mem_stage_inst_dmem_ram_177__3_), .D(
        mem_stage_inst_dmem_ram_179__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n499) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u934 ( .A(
        mem_stage_inst_dmem_ram_144__3_), .B(mem_stage_inst_dmem_ram_146__3_), 
        .C(mem_stage_inst_dmem_ram_145__3_), .D(
        mem_stage_inst_dmem_ram_147__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n509) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u933 ( .A(
        mem_stage_inst_dmem_ram_128__3_), .B(mem_stage_inst_dmem_ram_130__3_), 
        .C(mem_stage_inst_dmem_ram_129__3_), .D(
        mem_stage_inst_dmem_ram_131__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n514) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u932 ( .A(mem_stage_inst_dmem_ram_48__2_), .B(mem_stage_inst_dmem_ram_50__2_), .C(mem_stage_inst_dmem_ram_49__2_), .D(
        mem_stage_inst_dmem_ram_51__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n455) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u931 ( .A(mem_stage_inst_dmem_ram_16__2_), .B(mem_stage_inst_dmem_ram_18__2_), .C(mem_stage_inst_dmem_ram_17__2_), .D(
        mem_stage_inst_dmem_ram_19__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n465) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u930 ( .A(mem_stage_inst_dmem_ram_0__2_), 
        .B(mem_stage_inst_dmem_ram_2__2_), .C(mem_stage_inst_dmem_ram_1__2_), 
        .D(mem_stage_inst_dmem_ram_3__2_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n470) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u929 ( .A(
        mem_stage_inst_dmem_ram_176__2_), .B(mem_stage_inst_dmem_ram_178__2_), 
        .C(mem_stage_inst_dmem_ram_177__2_), .D(
        mem_stage_inst_dmem_ram_179__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n415) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u928 ( .A(
        mem_stage_inst_dmem_ram_144__2_), .B(mem_stage_inst_dmem_ram_146__2_), 
        .C(mem_stage_inst_dmem_ram_145__2_), .D(
        mem_stage_inst_dmem_ram_147__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n425) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u927 ( .A(
        mem_stage_inst_dmem_ram_128__2_), .B(mem_stage_inst_dmem_ram_130__2_), 
        .C(mem_stage_inst_dmem_ram_129__2_), .D(
        mem_stage_inst_dmem_ram_131__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n430) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u926 ( .A(mem_stage_inst_dmem_ram_48__1_), .B(mem_stage_inst_dmem_ram_50__1_), .C(mem_stage_inst_dmem_ram_49__1_), .D(
        mem_stage_inst_dmem_ram_51__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n371) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u925 ( .A(mem_stage_inst_dmem_ram_16__1_), .B(mem_stage_inst_dmem_ram_18__1_), .C(mem_stage_inst_dmem_ram_17__1_), .D(
        mem_stage_inst_dmem_ram_19__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n381) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u924 ( .A(mem_stage_inst_dmem_ram_0__1_), 
        .B(mem_stage_inst_dmem_ram_2__1_), .C(mem_stage_inst_dmem_ram_1__1_), 
        .D(mem_stage_inst_dmem_ram_3__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n386) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u923 ( .A(
        mem_stage_inst_dmem_ram_176__1_), .B(mem_stage_inst_dmem_ram_178__1_), 
        .C(mem_stage_inst_dmem_ram_177__1_), .D(
        mem_stage_inst_dmem_ram_179__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n331) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u922 ( .A(
        mem_stage_inst_dmem_ram_144__1_), .B(mem_stage_inst_dmem_ram_146__1_), 
        .C(mem_stage_inst_dmem_ram_145__1_), .D(
        mem_stage_inst_dmem_ram_147__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n341) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u921 ( .A(
        mem_stage_inst_dmem_ram_128__1_), .B(mem_stage_inst_dmem_ram_130__1_), 
        .C(mem_stage_inst_dmem_ram_129__1_), .D(
        mem_stage_inst_dmem_ram_131__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n346) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u920 ( .A(mem_stage_inst_dmem_ram_48__0_), .B(mem_stage_inst_dmem_ram_50__0_), .C(mem_stage_inst_dmem_ram_49__0_), .D(
        mem_stage_inst_dmem_ram_51__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n287) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u919 ( .A(mem_stage_inst_dmem_ram_16__0_), .B(mem_stage_inst_dmem_ram_18__0_), .C(mem_stage_inst_dmem_ram_17__0_), .D(
        mem_stage_inst_dmem_ram_19__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n297) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u918 ( .A(mem_stage_inst_dmem_ram_0__0_), 
        .B(mem_stage_inst_dmem_ram_2__0_), .C(mem_stage_inst_dmem_ram_1__0_), 
        .D(mem_stage_inst_dmem_ram_3__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n302) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u917 ( .A(
        mem_stage_inst_dmem_ram_176__0_), .B(mem_stage_inst_dmem_ram_178__0_), 
        .C(mem_stage_inst_dmem_ram_177__0_), .D(
        mem_stage_inst_dmem_ram_179__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n247) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u916 ( .A(
        mem_stage_inst_dmem_ram_144__0_), .B(mem_stage_inst_dmem_ram_146__0_), 
        .C(mem_stage_inst_dmem_ram_145__0_), .D(
        mem_stage_inst_dmem_ram_147__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n257) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u915 ( .A(
        mem_stage_inst_dmem_ram_128__0_), .B(mem_stage_inst_dmem_ram_130__0_), 
        .C(mem_stage_inst_dmem_ram_129__0_), .D(
        mem_stage_inst_dmem_ram_131__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n262) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u914 ( .A(
        mem_stage_inst_dmem_ram_224__15_), .B(mem_stage_inst_dmem_ram_226__15_), .C(mem_stage_inst_dmem_ram_225__15_), .D(mem_stage_inst_dmem_ram_227__15_), 
        .S0(mem_stage_inst_dmem_n138), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5588) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u913 ( .A(
        mem_stage_inst_dmem_ram_228__15_), .B(mem_stage_inst_dmem_ram_230__15_), .C(mem_stage_inst_dmem_ram_229__15_), .D(mem_stage_inst_dmem_ram_231__15_), 
        .S0(mem_stage_inst_dmem_n137), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5590) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u912 ( .A(
        mem_stage_inst_dmem_ram_236__15_), .B(mem_stage_inst_dmem_ram_238__15_), .C(mem_stage_inst_dmem_ram_237__15_), .D(mem_stage_inst_dmem_ram_239__15_), 
        .S0(mem_stage_inst_dmem_n136), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5591) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u911 ( .A(mem_stage_inst_dmem_n5588), 
        .B(mem_stage_inst_dmem_n5589), .C(mem_stage_inst_dmem_n5590), .D(
        mem_stage_inst_dmem_n5591), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5587) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u910 ( .A(
        mem_stage_inst_dmem_ram_96__15_), .B(mem_stage_inst_dmem_ram_98__15_), 
        .C(mem_stage_inst_dmem_ram_97__15_), .D(
        mem_stage_inst_dmem_ram_99__15_), .S0(ex_pipeline_reg_out[23]), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n5628) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u909 ( .A(
        mem_stage_inst_dmem_ram_100__15_), .B(mem_stage_inst_dmem_ram_102__15_), .C(mem_stage_inst_dmem_ram_101__15_), .D(mem_stage_inst_dmem_ram_103__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n36), .Y(
        mem_stage_inst_dmem_n5630) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u908 ( .A(
        mem_stage_inst_dmem_ram_108__15_), .B(mem_stage_inst_dmem_ram_110__15_), .C(mem_stage_inst_dmem_ram_109__15_), .D(mem_stage_inst_dmem_ram_111__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n35), .Y(
        mem_stage_inst_dmem_n5631) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u907 ( .A(mem_stage_inst_dmem_n5628), 
        .B(mem_stage_inst_dmem_n5629), .C(mem_stage_inst_dmem_n5630), .D(
        mem_stage_inst_dmem_n5631), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5627) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u906 ( .A(
        mem_stage_inst_dmem_ram_32__15_), .B(mem_stage_inst_dmem_ram_34__15_), 
        .C(mem_stage_inst_dmem_ram_33__15_), .D(
        mem_stage_inst_dmem_ram_35__15_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n25), .Y(mem_stage_inst_dmem_n5648) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u905 ( .A(
        mem_stage_inst_dmem_ram_36__15_), .B(mem_stage_inst_dmem_ram_38__15_), 
        .C(mem_stage_inst_dmem_ram_37__15_), .D(
        mem_stage_inst_dmem_ram_39__15_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n5650) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u904 ( .A(
        mem_stage_inst_dmem_ram_44__15_), .B(mem_stage_inst_dmem_ram_46__15_), 
        .C(mem_stage_inst_dmem_ram_45__15_), .D(
        mem_stage_inst_dmem_ram_47__15_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n5651) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u903 ( .A(mem_stage_inst_dmem_n5648), 
        .B(mem_stage_inst_dmem_n5649), .C(mem_stage_inst_dmem_n5650), .D(
        mem_stage_inst_dmem_n5651), .S0(mem_stage_inst_dmem_n209), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5647) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u902 ( .A(
        mem_stage_inst_dmem_ram_160__15_), .B(mem_stage_inst_dmem_ram_162__15_), .C(mem_stage_inst_dmem_ram_161__15_), .D(mem_stage_inst_dmem_ram_163__15_), 
        .S0(mem_stage_inst_dmem_n163), .S1(mem_stage_inst_dmem_n17), .Y(
        mem_stage_inst_dmem_n5608) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u901 ( .A(
        mem_stage_inst_dmem_ram_164__15_), .B(mem_stage_inst_dmem_ram_166__15_), .C(mem_stage_inst_dmem_ram_165__15_), .D(mem_stage_inst_dmem_ram_167__15_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n18), .Y(
        mem_stage_inst_dmem_n5610) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u900 ( .A(
        mem_stage_inst_dmem_ram_172__15_), .B(mem_stage_inst_dmem_ram_174__15_), .C(mem_stage_inst_dmem_ram_173__15_), .D(mem_stage_inst_dmem_ram_175__15_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n15), .Y(
        mem_stage_inst_dmem_n5611) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u899 ( .A(mem_stage_inst_dmem_n5608), 
        .B(mem_stage_inst_dmem_n5609), .C(mem_stage_inst_dmem_n5610), .D(
        mem_stage_inst_dmem_n5611), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5607) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u898 ( .A(
        mem_stage_inst_dmem_ram_224__14_), .B(mem_stage_inst_dmem_ram_226__14_), .C(mem_stage_inst_dmem_ram_225__14_), .D(mem_stage_inst_dmem_ram_227__14_), 
        .S0(mem_stage_inst_dmem_n120), .S1(mem_stage_inst_dmem_n56), .Y(
        mem_stage_inst_dmem_n5504) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u897 ( .A(
        mem_stage_inst_dmem_ram_228__14_), .B(mem_stage_inst_dmem_ram_230__14_), .C(mem_stage_inst_dmem_ram_229__14_), .D(mem_stage_inst_dmem_ram_231__14_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n55), .Y(
        mem_stage_inst_dmem_n5506) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u896 ( .A(
        mem_stage_inst_dmem_ram_236__14_), .B(mem_stage_inst_dmem_ram_238__14_), .C(mem_stage_inst_dmem_ram_237__14_), .D(mem_stage_inst_dmem_ram_239__14_), 
        .S0(mem_stage_inst_dmem_n108), .S1(mem_stage_inst_dmem_n54), .Y(
        mem_stage_inst_dmem_n5507) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u895 ( .A(mem_stage_inst_dmem_n5504), 
        .B(mem_stage_inst_dmem_n5505), .C(mem_stage_inst_dmem_n5506), .D(
        mem_stage_inst_dmem_n5507), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5503) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u894 ( .A(
        mem_stage_inst_dmem_ram_96__14_), .B(mem_stage_inst_dmem_ram_98__14_), 
        .C(mem_stage_inst_dmem_ram_97__14_), .D(
        mem_stage_inst_dmem_ram_99__14_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5544) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u893 ( .A(
        mem_stage_inst_dmem_ram_100__14_), .B(mem_stage_inst_dmem_ram_102__14_), .C(mem_stage_inst_dmem_ram_101__14_), .D(mem_stage_inst_dmem_ram_103__14_), 
        .S0(mem_stage_inst_dmem_n151), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5546) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u892 ( .A(
        mem_stage_inst_dmem_ram_108__14_), .B(mem_stage_inst_dmem_ram_110__14_), .C(mem_stage_inst_dmem_ram_109__14_), .D(mem_stage_inst_dmem_ram_111__14_), 
        .S0(mem_stage_inst_dmem_n149), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5547) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u891 ( .A(mem_stage_inst_dmem_n5544), 
        .B(mem_stage_inst_dmem_n5545), .C(mem_stage_inst_dmem_n5546), .D(
        mem_stage_inst_dmem_n5547), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5543) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u890 ( .A(
        mem_stage_inst_dmem_ram_32__14_), .B(mem_stage_inst_dmem_ram_34__14_), 
        .C(mem_stage_inst_dmem_ram_33__14_), .D(
        mem_stage_inst_dmem_ram_35__14_), .S0(mem_stage_inst_dmem_n117), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5564) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u889 ( .A(
        mem_stage_inst_dmem_ram_36__14_), .B(mem_stage_inst_dmem_ram_38__14_), 
        .C(mem_stage_inst_dmem_ram_37__14_), .D(
        mem_stage_inst_dmem_ram_39__14_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5566) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u888 ( .A(
        mem_stage_inst_dmem_ram_44__14_), .B(mem_stage_inst_dmem_ram_46__14_), 
        .C(mem_stage_inst_dmem_ram_45__14_), .D(
        mem_stage_inst_dmem_ram_47__14_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5567) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u887 ( .A(mem_stage_inst_dmem_n5564), 
        .B(mem_stage_inst_dmem_n5565), .C(mem_stage_inst_dmem_n5566), .D(
        mem_stage_inst_dmem_n5567), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5563) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u886 ( .A(
        mem_stage_inst_dmem_ram_160__14_), .B(mem_stage_inst_dmem_ram_162__14_), .C(mem_stage_inst_dmem_ram_161__14_), .D(mem_stage_inst_dmem_ram_163__14_), 
        .S0(mem_stage_inst_dmem_n164), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5524) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u885 ( .A(
        mem_stage_inst_dmem_ram_164__14_), .B(mem_stage_inst_dmem_ram_166__14_), .C(mem_stage_inst_dmem_ram_165__14_), .D(mem_stage_inst_dmem_ram_167__14_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5526) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u884 ( .A(
        mem_stage_inst_dmem_ram_172__14_), .B(mem_stage_inst_dmem_ram_174__14_), .C(mem_stage_inst_dmem_ram_173__14_), .D(mem_stage_inst_dmem_ram_175__14_), 
        .S0(mem_stage_inst_dmem_n110), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5527) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u883 ( .A(mem_stage_inst_dmem_n5524), 
        .B(mem_stage_inst_dmem_n5525), .C(mem_stage_inst_dmem_n5526), .D(
        mem_stage_inst_dmem_n5527), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5523) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u882 ( .A(
        mem_stage_inst_dmem_ram_224__13_), .B(mem_stage_inst_dmem_ram_226__13_), .C(mem_stage_inst_dmem_ram_225__13_), .D(mem_stage_inst_dmem_ram_227__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n37), .Y(
        mem_stage_inst_dmem_n5420) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u881 ( .A(
        mem_stage_inst_dmem_ram_228__13_), .B(mem_stage_inst_dmem_ram_230__13_), .C(mem_stage_inst_dmem_ram_229__13_), .D(mem_stage_inst_dmem_ram_231__13_), 
        .S0(mem_stage_inst_dmem_n147), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5422) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u880 ( .A(
        mem_stage_inst_dmem_ram_236__13_), .B(mem_stage_inst_dmem_ram_238__13_), .C(mem_stage_inst_dmem_ram_237__13_), .D(mem_stage_inst_dmem_ram_239__13_), 
        .S0(mem_stage_inst_dmem_n146), .S1(mem_stage_inst_dmem_n64), .Y(
        mem_stage_inst_dmem_n5423) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u879 ( .A(mem_stage_inst_dmem_n5420), 
        .B(mem_stage_inst_dmem_n5421), .C(mem_stage_inst_dmem_n5422), .D(
        mem_stage_inst_dmem_n5423), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5419) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u878 ( .A(
        mem_stage_inst_dmem_ram_96__13_), .B(mem_stage_inst_dmem_ram_98__13_), 
        .C(mem_stage_inst_dmem_ram_97__13_), .D(
        mem_stage_inst_dmem_ram_99__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n5460) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u877 ( .A(
        mem_stage_inst_dmem_ram_100__13_), .B(mem_stage_inst_dmem_ram_102__13_), .C(mem_stage_inst_dmem_ram_101__13_), .D(mem_stage_inst_dmem_ram_103__13_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n60), .Y(
        mem_stage_inst_dmem_n5462) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u876 ( .A(
        mem_stage_inst_dmem_ram_108__13_), .B(mem_stage_inst_dmem_ram_110__13_), .C(mem_stage_inst_dmem_ram_109__13_), .D(mem_stage_inst_dmem_ram_111__13_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n59), .Y(
        mem_stage_inst_dmem_n5463) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u875 ( .A(mem_stage_inst_dmem_n5460), 
        .B(mem_stage_inst_dmem_n5461), .C(mem_stage_inst_dmem_n5462), .D(
        mem_stage_inst_dmem_n5463), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5459) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u874 ( .A(
        mem_stage_inst_dmem_ram_32__13_), .B(mem_stage_inst_dmem_ram_34__13_), 
        .C(mem_stage_inst_dmem_ram_33__13_), .D(
        mem_stage_inst_dmem_ram_35__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5480) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u873 ( .A(
        mem_stage_inst_dmem_ram_36__13_), .B(mem_stage_inst_dmem_ram_38__13_), 
        .C(mem_stage_inst_dmem_ram_37__13_), .D(
        mem_stage_inst_dmem_ram_39__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5482) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u872 ( .A(
        mem_stage_inst_dmem_ram_44__13_), .B(mem_stage_inst_dmem_ram_46__13_), 
        .C(mem_stage_inst_dmem_ram_45__13_), .D(
        mem_stage_inst_dmem_ram_47__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5483) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u871 ( .A(mem_stage_inst_dmem_n5480), 
        .B(mem_stage_inst_dmem_n5481), .C(mem_stage_inst_dmem_n5482), .D(
        mem_stage_inst_dmem_n5483), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5479) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u870 ( .A(
        mem_stage_inst_dmem_ram_160__13_), .B(mem_stage_inst_dmem_ram_162__13_), .C(mem_stage_inst_dmem_ram_161__13_), .D(mem_stage_inst_dmem_ram_163__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5440) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u869 ( .A(
        mem_stage_inst_dmem_ram_164__13_), .B(mem_stage_inst_dmem_ram_166__13_), .C(mem_stage_inst_dmem_ram_165__13_), .D(mem_stage_inst_dmem_ram_167__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5442) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u868 ( .A(
        mem_stage_inst_dmem_ram_172__13_), .B(mem_stage_inst_dmem_ram_174__13_), .C(mem_stage_inst_dmem_ram_173__13_), .D(mem_stage_inst_dmem_ram_175__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5443) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u867 ( .A(mem_stage_inst_dmem_n5440), 
        .B(mem_stage_inst_dmem_n5441), .C(mem_stage_inst_dmem_n5442), .D(
        mem_stage_inst_dmem_n5443), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5439) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u866 ( .A(
        mem_stage_inst_dmem_ram_224__12_), .B(mem_stage_inst_dmem_ram_226__12_), .C(mem_stage_inst_dmem_ram_225__12_), .D(mem_stage_inst_dmem_ram_227__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5336) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u865 ( .A(
        mem_stage_inst_dmem_ram_228__12_), .B(mem_stage_inst_dmem_ram_230__12_), .C(mem_stage_inst_dmem_ram_229__12_), .D(mem_stage_inst_dmem_ram_231__12_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n47), .Y(
        mem_stage_inst_dmem_n5338) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u864 ( .A(
        mem_stage_inst_dmem_ram_236__12_), .B(mem_stage_inst_dmem_ram_238__12_), .C(mem_stage_inst_dmem_ram_237__12_), .D(mem_stage_inst_dmem_ram_239__12_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n27), .Y(
        mem_stage_inst_dmem_n5339) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u863 ( .A(mem_stage_inst_dmem_n5336), 
        .B(mem_stage_inst_dmem_n5337), .C(mem_stage_inst_dmem_n5338), .D(
        mem_stage_inst_dmem_n5339), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5335) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u862 ( .A(
        mem_stage_inst_dmem_ram_96__12_), .B(mem_stage_inst_dmem_ram_98__12_), 
        .C(mem_stage_inst_dmem_ram_97__12_), .D(
        mem_stage_inst_dmem_ram_99__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5376) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u861 ( .A(
        mem_stage_inst_dmem_ram_100__12_), .B(mem_stage_inst_dmem_ram_102__12_), .C(mem_stage_inst_dmem_ram_101__12_), .D(mem_stage_inst_dmem_ram_103__12_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5378) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u860 ( .A(
        mem_stage_inst_dmem_ram_108__12_), .B(mem_stage_inst_dmem_ram_110__12_), .C(mem_stage_inst_dmem_ram_109__12_), .D(mem_stage_inst_dmem_ram_111__12_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5379) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u859 ( .A(mem_stage_inst_dmem_n5376), 
        .B(mem_stage_inst_dmem_n5377), .C(mem_stage_inst_dmem_n5378), .D(
        mem_stage_inst_dmem_n5379), .S0(mem_stage_inst_dmem_n217), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5375) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u858 ( .A(
        mem_stage_inst_dmem_ram_32__12_), .B(mem_stage_inst_dmem_ram_34__12_), 
        .C(mem_stage_inst_dmem_ram_33__12_), .D(
        mem_stage_inst_dmem_ram_35__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n5396) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u857 ( .A(
        mem_stage_inst_dmem_ram_36__12_), .B(mem_stage_inst_dmem_ram_38__12_), 
        .C(mem_stage_inst_dmem_ram_37__12_), .D(
        mem_stage_inst_dmem_ram_39__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n5398) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u856 ( .A(
        mem_stage_inst_dmem_ram_44__12_), .B(mem_stage_inst_dmem_ram_46__12_), 
        .C(mem_stage_inst_dmem_ram_45__12_), .D(
        mem_stage_inst_dmem_ram_47__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n5399) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u855 ( .A(mem_stage_inst_dmem_n5396), 
        .B(mem_stage_inst_dmem_n5397), .C(mem_stage_inst_dmem_n5398), .D(
        mem_stage_inst_dmem_n5399), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5395) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u854 ( .A(
        mem_stage_inst_dmem_ram_160__12_), .B(mem_stage_inst_dmem_ram_162__12_), .C(mem_stage_inst_dmem_ram_161__12_), .D(mem_stage_inst_dmem_ram_163__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5356) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u853 ( .A(
        mem_stage_inst_dmem_ram_164__12_), .B(mem_stage_inst_dmem_ram_166__12_), .C(mem_stage_inst_dmem_ram_165__12_), .D(mem_stage_inst_dmem_ram_167__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5358) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u852 ( .A(
        mem_stage_inst_dmem_ram_172__12_), .B(mem_stage_inst_dmem_ram_174__12_), .C(mem_stage_inst_dmem_ram_173__12_), .D(mem_stage_inst_dmem_ram_175__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5359) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u851 ( .A(mem_stage_inst_dmem_n5356), 
        .B(mem_stage_inst_dmem_n5357), .C(mem_stage_inst_dmem_n5358), .D(
        mem_stage_inst_dmem_n5359), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5355) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u850 ( .A(
        mem_stage_inst_dmem_ram_224__11_), .B(mem_stage_inst_dmem_ram_226__11_), .C(mem_stage_inst_dmem_ram_225__11_), .D(mem_stage_inst_dmem_ram_227__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5252) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u849 ( .A(
        mem_stage_inst_dmem_ram_228__11_), .B(mem_stage_inst_dmem_ram_230__11_), .C(mem_stage_inst_dmem_ram_229__11_), .D(mem_stage_inst_dmem_ram_231__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5254) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u848 ( .A(
        mem_stage_inst_dmem_ram_236__11_), .B(mem_stage_inst_dmem_ram_238__11_), .C(mem_stage_inst_dmem_ram_237__11_), .D(mem_stage_inst_dmem_ram_239__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5255) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u847 ( .A(mem_stage_inst_dmem_n5252), 
        .B(mem_stage_inst_dmem_n5253), .C(mem_stage_inst_dmem_n5254), .D(
        mem_stage_inst_dmem_n5255), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5251) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u846 ( .A(
        mem_stage_inst_dmem_ram_96__11_), .B(mem_stage_inst_dmem_ram_98__11_), 
        .C(mem_stage_inst_dmem_ram_97__11_), .D(
        mem_stage_inst_dmem_ram_99__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5292) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u845 ( .A(
        mem_stage_inst_dmem_ram_100__11_), .B(mem_stage_inst_dmem_ram_102__11_), .C(mem_stage_inst_dmem_ram_101__11_), .D(mem_stage_inst_dmem_ram_103__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5294) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u844 ( .A(
        mem_stage_inst_dmem_ram_108__11_), .B(mem_stage_inst_dmem_ram_110__11_), .C(mem_stage_inst_dmem_ram_109__11_), .D(mem_stage_inst_dmem_ram_111__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5295) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u843 ( .A(mem_stage_inst_dmem_n5292), 
        .B(mem_stage_inst_dmem_n5293), .C(mem_stage_inst_dmem_n5294), .D(
        mem_stage_inst_dmem_n5295), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5291) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u842 ( .A(
        mem_stage_inst_dmem_ram_32__11_), .B(mem_stage_inst_dmem_ram_34__11_), 
        .C(mem_stage_inst_dmem_ram_33__11_), .D(
        mem_stage_inst_dmem_ram_35__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5312) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u841 ( .A(
        mem_stage_inst_dmem_ram_36__11_), .B(mem_stage_inst_dmem_ram_38__11_), 
        .C(mem_stage_inst_dmem_ram_37__11_), .D(
        mem_stage_inst_dmem_ram_39__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5314) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u840 ( .A(
        mem_stage_inst_dmem_ram_44__11_), .B(mem_stage_inst_dmem_ram_46__11_), 
        .C(mem_stage_inst_dmem_ram_45__11_), .D(
        mem_stage_inst_dmem_ram_47__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5315) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u839 ( .A(mem_stage_inst_dmem_n5312), 
        .B(mem_stage_inst_dmem_n5313), .C(mem_stage_inst_dmem_n5314), .D(
        mem_stage_inst_dmem_n5315), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5311) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u838 ( .A(
        mem_stage_inst_dmem_ram_160__11_), .B(mem_stage_inst_dmem_ram_162__11_), .C(mem_stage_inst_dmem_ram_161__11_), .D(mem_stage_inst_dmem_ram_163__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5272) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u837 ( .A(
        mem_stage_inst_dmem_ram_164__11_), .B(mem_stage_inst_dmem_ram_166__11_), .C(mem_stage_inst_dmem_ram_165__11_), .D(mem_stage_inst_dmem_ram_167__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5274) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u836 ( .A(
        mem_stage_inst_dmem_ram_172__11_), .B(mem_stage_inst_dmem_ram_174__11_), .C(mem_stage_inst_dmem_ram_173__11_), .D(mem_stage_inst_dmem_ram_175__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5275) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u835 ( .A(mem_stage_inst_dmem_n5272), 
        .B(mem_stage_inst_dmem_n5273), .C(mem_stage_inst_dmem_n5274), .D(
        mem_stage_inst_dmem_n5275), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5271) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u834 ( .A(
        mem_stage_inst_dmem_ram_224__10_), .B(mem_stage_inst_dmem_ram_226__10_), .C(mem_stage_inst_dmem_ram_225__10_), .D(mem_stage_inst_dmem_ram_227__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5168) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u833 ( .A(
        mem_stage_inst_dmem_ram_228__10_), .B(mem_stage_inst_dmem_ram_230__10_), .C(mem_stage_inst_dmem_ram_229__10_), .D(mem_stage_inst_dmem_ram_231__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5170) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u832 ( .A(
        mem_stage_inst_dmem_ram_236__10_), .B(mem_stage_inst_dmem_ram_238__10_), .C(mem_stage_inst_dmem_ram_237__10_), .D(mem_stage_inst_dmem_ram_239__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5171) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u831 ( .A(mem_stage_inst_dmem_n5168), 
        .B(mem_stage_inst_dmem_n5169), .C(mem_stage_inst_dmem_n5170), .D(
        mem_stage_inst_dmem_n5171), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5167) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u830 ( .A(
        mem_stage_inst_dmem_ram_96__10_), .B(mem_stage_inst_dmem_ram_98__10_), 
        .C(mem_stage_inst_dmem_ram_97__10_), .D(
        mem_stage_inst_dmem_ram_99__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5208) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u829 ( .A(
        mem_stage_inst_dmem_ram_100__10_), .B(mem_stage_inst_dmem_ram_102__10_), .C(mem_stage_inst_dmem_ram_101__10_), .D(mem_stage_inst_dmem_ram_103__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5210) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u828 ( .A(
        mem_stage_inst_dmem_ram_108__10_), .B(mem_stage_inst_dmem_ram_110__10_), .C(mem_stage_inst_dmem_ram_109__10_), .D(mem_stage_inst_dmem_ram_111__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5211) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u827 ( .A(mem_stage_inst_dmem_n5208), 
        .B(mem_stage_inst_dmem_n5209), .C(mem_stage_inst_dmem_n5210), .D(
        mem_stage_inst_dmem_n5211), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5207) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u826 ( .A(
        mem_stage_inst_dmem_ram_32__10_), .B(mem_stage_inst_dmem_ram_34__10_), 
        .C(mem_stage_inst_dmem_ram_33__10_), .D(
        mem_stage_inst_dmem_ram_35__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5228) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u825 ( .A(
        mem_stage_inst_dmem_ram_36__10_), .B(mem_stage_inst_dmem_ram_38__10_), 
        .C(mem_stage_inst_dmem_ram_37__10_), .D(
        mem_stage_inst_dmem_ram_39__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5230) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u824 ( .A(
        mem_stage_inst_dmem_ram_44__10_), .B(mem_stage_inst_dmem_ram_46__10_), 
        .C(mem_stage_inst_dmem_ram_45__10_), .D(
        mem_stage_inst_dmem_ram_47__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5231) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u823 ( .A(mem_stage_inst_dmem_n5228), 
        .B(mem_stage_inst_dmem_n5229), .C(mem_stage_inst_dmem_n5230), .D(
        mem_stage_inst_dmem_n5231), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5227) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u822 ( .A(
        mem_stage_inst_dmem_ram_160__10_), .B(mem_stage_inst_dmem_ram_162__10_), .C(mem_stage_inst_dmem_ram_161__10_), .D(mem_stage_inst_dmem_ram_163__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5188) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u821 ( .A(
        mem_stage_inst_dmem_ram_164__10_), .B(mem_stage_inst_dmem_ram_166__10_), .C(mem_stage_inst_dmem_ram_165__10_), .D(mem_stage_inst_dmem_ram_167__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5190) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u820 ( .A(
        mem_stage_inst_dmem_ram_172__10_), .B(mem_stage_inst_dmem_ram_174__10_), .C(mem_stage_inst_dmem_ram_173__10_), .D(mem_stage_inst_dmem_ram_175__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5191) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u819 ( .A(mem_stage_inst_dmem_n5188), 
        .B(mem_stage_inst_dmem_n5189), .C(mem_stage_inst_dmem_n5190), .D(
        mem_stage_inst_dmem_n5191), .S0(ex_pipeline_reg_out[25]), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5187) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u818 ( .A(
        mem_stage_inst_dmem_ram_224__9_), .B(mem_stage_inst_dmem_ram_226__9_), 
        .C(mem_stage_inst_dmem_ram_225__9_), .D(
        mem_stage_inst_dmem_ram_227__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5084) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u817 ( .A(
        mem_stage_inst_dmem_ram_228__9_), .B(mem_stage_inst_dmem_ram_230__9_), 
        .C(mem_stage_inst_dmem_ram_229__9_), .D(
        mem_stage_inst_dmem_ram_231__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5086) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u816 ( .A(
        mem_stage_inst_dmem_ram_236__9_), .B(mem_stage_inst_dmem_ram_238__9_), 
        .C(mem_stage_inst_dmem_ram_237__9_), .D(
        mem_stage_inst_dmem_ram_239__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5087) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u815 ( .A(mem_stage_inst_dmem_n5084), 
        .B(mem_stage_inst_dmem_n5085), .C(mem_stage_inst_dmem_n5086), .D(
        mem_stage_inst_dmem_n5087), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5083) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u814 ( .A(mem_stage_inst_dmem_ram_96__9_), .B(mem_stage_inst_dmem_ram_98__9_), .C(mem_stage_inst_dmem_ram_97__9_), .D(
        mem_stage_inst_dmem_ram_99__9_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5124) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u813 ( .A(
        mem_stage_inst_dmem_ram_100__9_), .B(mem_stage_inst_dmem_ram_102__9_), 
        .C(mem_stage_inst_dmem_ram_101__9_), .D(
        mem_stage_inst_dmem_ram_103__9_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5126) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u812 ( .A(
        mem_stage_inst_dmem_ram_108__9_), .B(mem_stage_inst_dmem_ram_110__9_), 
        .C(mem_stage_inst_dmem_ram_109__9_), .D(
        mem_stage_inst_dmem_ram_111__9_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5127) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u811 ( .A(mem_stage_inst_dmem_n5124), 
        .B(mem_stage_inst_dmem_n5125), .C(mem_stage_inst_dmem_n5126), .D(
        mem_stage_inst_dmem_n5127), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5123) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u810 ( .A(mem_stage_inst_dmem_ram_32__9_), .B(mem_stage_inst_dmem_ram_34__9_), .C(mem_stage_inst_dmem_ram_33__9_), .D(
        mem_stage_inst_dmem_ram_35__9_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n5144) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u809 ( .A(mem_stage_inst_dmem_ram_36__9_), .B(mem_stage_inst_dmem_ram_38__9_), .C(mem_stage_inst_dmem_ram_37__9_), .D(
        mem_stage_inst_dmem_ram_39__9_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n19), .Y(mem_stage_inst_dmem_n5146) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u808 ( .A(mem_stage_inst_dmem_ram_44__9_), .B(mem_stage_inst_dmem_ram_46__9_), .C(mem_stage_inst_dmem_ram_45__9_), .D(
        mem_stage_inst_dmem_ram_47__9_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5147) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u807 ( .A(mem_stage_inst_dmem_n5144), 
        .B(mem_stage_inst_dmem_n5145), .C(mem_stage_inst_dmem_n5146), .D(
        mem_stage_inst_dmem_n5147), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5143) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u806 ( .A(
        mem_stage_inst_dmem_ram_160__9_), .B(mem_stage_inst_dmem_ram_162__9_), 
        .C(mem_stage_inst_dmem_ram_161__9_), .D(
        mem_stage_inst_dmem_ram_163__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5104) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u805 ( .A(
        mem_stage_inst_dmem_ram_164__9_), .B(mem_stage_inst_dmem_ram_166__9_), 
        .C(mem_stage_inst_dmem_ram_165__9_), .D(
        mem_stage_inst_dmem_ram_167__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5106) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u804 ( .A(
        mem_stage_inst_dmem_ram_172__9_), .B(mem_stage_inst_dmem_ram_174__9_), 
        .C(mem_stage_inst_dmem_ram_173__9_), .D(
        mem_stage_inst_dmem_ram_175__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5107) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u803 ( .A(mem_stage_inst_dmem_n5104), 
        .B(mem_stage_inst_dmem_n5105), .C(mem_stage_inst_dmem_n5106), .D(
        mem_stage_inst_dmem_n5107), .S0(mem_stage_inst_dmem_n214), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5103) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u802 ( .A(
        mem_stage_inst_dmem_ram_224__8_), .B(mem_stage_inst_dmem_ram_226__8_), 
        .C(mem_stage_inst_dmem_ram_225__8_), .D(
        mem_stage_inst_dmem_ram_227__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5000) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u801 ( .A(
        mem_stage_inst_dmem_ram_228__8_), .B(mem_stage_inst_dmem_ram_230__8_), 
        .C(mem_stage_inst_dmem_ram_229__8_), .D(
        mem_stage_inst_dmem_ram_231__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5002) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u800 ( .A(
        mem_stage_inst_dmem_ram_236__8_), .B(mem_stage_inst_dmem_ram_238__8_), 
        .C(mem_stage_inst_dmem_ram_237__8_), .D(
        mem_stage_inst_dmem_ram_239__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5003) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u799 ( .A(mem_stage_inst_dmem_n5000), 
        .B(mem_stage_inst_dmem_n5001), .C(mem_stage_inst_dmem_n5002), .D(
        mem_stage_inst_dmem_n5003), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4999) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u798 ( .A(mem_stage_inst_dmem_ram_96__8_), .B(mem_stage_inst_dmem_ram_98__8_), .C(mem_stage_inst_dmem_ram_97__8_), .D(
        mem_stage_inst_dmem_ram_99__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5040) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u797 ( .A(
        mem_stage_inst_dmem_ram_100__8_), .B(mem_stage_inst_dmem_ram_102__8_), 
        .C(mem_stage_inst_dmem_ram_101__8_), .D(
        mem_stage_inst_dmem_ram_103__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5042) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u796 ( .A(
        mem_stage_inst_dmem_ram_108__8_), .B(mem_stage_inst_dmem_ram_110__8_), 
        .C(mem_stage_inst_dmem_ram_109__8_), .D(
        mem_stage_inst_dmem_ram_111__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5043) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u795 ( .A(mem_stage_inst_dmem_n5040), 
        .B(mem_stage_inst_dmem_n5041), .C(mem_stage_inst_dmem_n5042), .D(
        mem_stage_inst_dmem_n5043), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5039) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u794 ( .A(mem_stage_inst_dmem_ram_32__8_), .B(mem_stage_inst_dmem_ram_34__8_), .C(mem_stage_inst_dmem_ram_33__8_), .D(
        mem_stage_inst_dmem_ram_35__8_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5060) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u793 ( .A(mem_stage_inst_dmem_ram_36__8_), .B(mem_stage_inst_dmem_ram_38__8_), .C(mem_stage_inst_dmem_ram_37__8_), .D(
        mem_stage_inst_dmem_ram_39__8_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5062) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u792 ( .A(mem_stage_inst_dmem_ram_44__8_), .B(mem_stage_inst_dmem_ram_46__8_), .C(mem_stage_inst_dmem_ram_45__8_), .D(
        mem_stage_inst_dmem_ram_47__8_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5063) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u791 ( .A(mem_stage_inst_dmem_n5060), 
        .B(mem_stage_inst_dmem_n5061), .C(mem_stage_inst_dmem_n5062), .D(
        mem_stage_inst_dmem_n5063), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5059) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u790 ( .A(
        mem_stage_inst_dmem_ram_160__8_), .B(mem_stage_inst_dmem_ram_162__8_), 
        .C(mem_stage_inst_dmem_ram_161__8_), .D(
        mem_stage_inst_dmem_ram_163__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5020) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u789 ( .A(
        mem_stage_inst_dmem_ram_164__8_), .B(mem_stage_inst_dmem_ram_166__8_), 
        .C(mem_stage_inst_dmem_ram_165__8_), .D(
        mem_stage_inst_dmem_ram_167__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5022) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u788 ( .A(
        mem_stage_inst_dmem_ram_172__8_), .B(mem_stage_inst_dmem_ram_174__8_), 
        .C(mem_stage_inst_dmem_ram_173__8_), .D(
        mem_stage_inst_dmem_ram_175__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5023) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u787 ( .A(mem_stage_inst_dmem_n5020), 
        .B(mem_stage_inst_dmem_n5021), .C(mem_stage_inst_dmem_n5022), .D(
        mem_stage_inst_dmem_n5023), .S0(mem_stage_inst_dmem_n213), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5019) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u786 ( .A(
        mem_stage_inst_dmem_ram_224__7_), .B(mem_stage_inst_dmem_ram_226__7_), 
        .C(mem_stage_inst_dmem_ram_225__7_), .D(
        mem_stage_inst_dmem_ram_227__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4916) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u785 ( .A(
        mem_stage_inst_dmem_ram_228__7_), .B(mem_stage_inst_dmem_ram_230__7_), 
        .C(mem_stage_inst_dmem_ram_229__7_), .D(
        mem_stage_inst_dmem_ram_231__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4918) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u784 ( .A(
        mem_stage_inst_dmem_ram_236__7_), .B(mem_stage_inst_dmem_ram_238__7_), 
        .C(mem_stage_inst_dmem_ram_237__7_), .D(
        mem_stage_inst_dmem_ram_239__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4919) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u783 ( .A(mem_stage_inst_dmem_n4916), 
        .B(mem_stage_inst_dmem_n4917), .C(mem_stage_inst_dmem_n4918), .D(
        mem_stage_inst_dmem_n4919), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4915) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u782 ( .A(mem_stage_inst_dmem_ram_96__7_), .B(mem_stage_inst_dmem_ram_98__7_), .C(mem_stage_inst_dmem_ram_97__7_), .D(
        mem_stage_inst_dmem_ram_99__7_), .S0(mem_stage_inst_dmem_n153), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n4956) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u781 ( .A(
        mem_stage_inst_dmem_ram_100__7_), .B(mem_stage_inst_dmem_ram_102__7_), 
        .C(mem_stage_inst_dmem_ram_101__7_), .D(
        mem_stage_inst_dmem_ram_103__7_), .S0(mem_stage_inst_dmem_n153), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n4958) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u780 ( .A(
        mem_stage_inst_dmem_ram_108__7_), .B(mem_stage_inst_dmem_ram_110__7_), 
        .C(mem_stage_inst_dmem_ram_109__7_), .D(
        mem_stage_inst_dmem_ram_111__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4959) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u779 ( .A(mem_stage_inst_dmem_n4956), 
        .B(mem_stage_inst_dmem_n4957), .C(mem_stage_inst_dmem_n4958), .D(
        mem_stage_inst_dmem_n4959), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4955) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u778 ( .A(mem_stage_inst_dmem_ram_32__7_), .B(mem_stage_inst_dmem_ram_34__7_), .C(mem_stage_inst_dmem_ram_33__7_), .D(
        mem_stage_inst_dmem_ram_35__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4976) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u777 ( .A(mem_stage_inst_dmem_ram_36__7_), .B(mem_stage_inst_dmem_ram_38__7_), .C(mem_stage_inst_dmem_ram_37__7_), .D(
        mem_stage_inst_dmem_ram_39__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4978) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u776 ( .A(mem_stage_inst_dmem_ram_44__7_), .B(mem_stage_inst_dmem_ram_46__7_), .C(mem_stage_inst_dmem_ram_45__7_), .D(
        mem_stage_inst_dmem_ram_47__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4979) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u775 ( .A(mem_stage_inst_dmem_n4976), 
        .B(mem_stage_inst_dmem_n4977), .C(mem_stage_inst_dmem_n4978), .D(
        mem_stage_inst_dmem_n4979), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4975) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u774 ( .A(
        mem_stage_inst_dmem_ram_160__7_), .B(mem_stage_inst_dmem_ram_162__7_), 
        .C(mem_stage_inst_dmem_ram_161__7_), .D(
        mem_stage_inst_dmem_ram_163__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4936) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u773 ( .A(
        mem_stage_inst_dmem_ram_164__7_), .B(mem_stage_inst_dmem_ram_166__7_), 
        .C(mem_stage_inst_dmem_ram_165__7_), .D(
        mem_stage_inst_dmem_ram_167__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4938) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u772 ( .A(
        mem_stage_inst_dmem_ram_172__7_), .B(mem_stage_inst_dmem_ram_174__7_), 
        .C(mem_stage_inst_dmem_ram_173__7_), .D(
        mem_stage_inst_dmem_ram_175__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4939) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u771 ( .A(mem_stage_inst_dmem_n4936), 
        .B(mem_stage_inst_dmem_n4937), .C(mem_stage_inst_dmem_n4938), .D(
        mem_stage_inst_dmem_n4939), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4935) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u770 ( .A(
        mem_stage_inst_dmem_ram_224__6_), .B(mem_stage_inst_dmem_ram_226__6_), 
        .C(mem_stage_inst_dmem_ram_225__6_), .D(
        mem_stage_inst_dmem_ram_227__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4832) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u769 ( .A(
        mem_stage_inst_dmem_ram_228__6_), .B(mem_stage_inst_dmem_ram_230__6_), 
        .C(mem_stage_inst_dmem_ram_229__6_), .D(
        mem_stage_inst_dmem_ram_231__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4834) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u768 ( .A(
        mem_stage_inst_dmem_ram_236__6_), .B(mem_stage_inst_dmem_ram_238__6_), 
        .C(mem_stage_inst_dmem_ram_237__6_), .D(
        mem_stage_inst_dmem_ram_239__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4835) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u767 ( .A(mem_stage_inst_dmem_n4832), 
        .B(mem_stage_inst_dmem_n4833), .C(mem_stage_inst_dmem_n4834), .D(
        mem_stage_inst_dmem_n4835), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4831) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u766 ( .A(mem_stage_inst_dmem_ram_96__6_), .B(mem_stage_inst_dmem_ram_98__6_), .C(mem_stage_inst_dmem_ram_97__6_), .D(
        mem_stage_inst_dmem_ram_99__6_), .S0(mem_stage_inst_dmem_n148), .S1(
        mem_stage_inst_dmem_n50), .Y(mem_stage_inst_dmem_n4872) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u765 ( .A(
        mem_stage_inst_dmem_ram_100__6_), .B(mem_stage_inst_dmem_ram_102__6_), 
        .C(mem_stage_inst_dmem_ram_101__6_), .D(
        mem_stage_inst_dmem_ram_103__6_), .S0(mem_stage_inst_dmem_n148), .S1(
        mem_stage_inst_dmem_n50), .Y(mem_stage_inst_dmem_n4874) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u764 ( .A(
        mem_stage_inst_dmem_ram_108__6_), .B(mem_stage_inst_dmem_ram_110__6_), 
        .C(mem_stage_inst_dmem_ram_109__6_), .D(
        mem_stage_inst_dmem_ram_111__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4875) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u763 ( .A(mem_stage_inst_dmem_n4872), 
        .B(mem_stage_inst_dmem_n4873), .C(mem_stage_inst_dmem_n4874), .D(
        mem_stage_inst_dmem_n4875), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4871) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u762 ( .A(mem_stage_inst_dmem_ram_32__6_), .B(mem_stage_inst_dmem_ram_34__6_), .C(mem_stage_inst_dmem_ram_33__6_), .D(
        mem_stage_inst_dmem_ram_35__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4892) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u761 ( .A(mem_stage_inst_dmem_ram_36__6_), .B(mem_stage_inst_dmem_ram_38__6_), .C(mem_stage_inst_dmem_ram_37__6_), .D(
        mem_stage_inst_dmem_ram_39__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4894) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u760 ( .A(mem_stage_inst_dmem_ram_44__6_), .B(mem_stage_inst_dmem_ram_46__6_), .C(mem_stage_inst_dmem_ram_45__6_), .D(
        mem_stage_inst_dmem_ram_47__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4895) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u759 ( .A(mem_stage_inst_dmem_n4892), 
        .B(mem_stage_inst_dmem_n4893), .C(mem_stage_inst_dmem_n4894), .D(
        mem_stage_inst_dmem_n4895), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4891) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u758 ( .A(
        mem_stage_inst_dmem_ram_160__6_), .B(mem_stage_inst_dmem_ram_162__6_), 
        .C(mem_stage_inst_dmem_ram_161__6_), .D(
        mem_stage_inst_dmem_ram_163__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4852) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u757 ( .A(
        mem_stage_inst_dmem_ram_164__6_), .B(mem_stage_inst_dmem_ram_166__6_), 
        .C(mem_stage_inst_dmem_ram_165__6_), .D(
        mem_stage_inst_dmem_ram_167__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4854) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u756 ( .A(
        mem_stage_inst_dmem_ram_172__6_), .B(mem_stage_inst_dmem_ram_174__6_), 
        .C(mem_stage_inst_dmem_ram_173__6_), .D(
        mem_stage_inst_dmem_ram_175__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4855) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u755 ( .A(mem_stage_inst_dmem_n4852), 
        .B(mem_stage_inst_dmem_n4853), .C(mem_stage_inst_dmem_n4854), .D(
        mem_stage_inst_dmem_n4855), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4851) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u754 ( .A(
        mem_stage_inst_dmem_ram_224__5_), .B(mem_stage_inst_dmem_ram_226__5_), 
        .C(mem_stage_inst_dmem_ram_225__5_), .D(
        mem_stage_inst_dmem_ram_227__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4748) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u753 ( .A(
        mem_stage_inst_dmem_ram_228__5_), .B(mem_stage_inst_dmem_ram_230__5_), 
        .C(mem_stage_inst_dmem_ram_229__5_), .D(
        mem_stage_inst_dmem_ram_231__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4750) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u752 ( .A(
        mem_stage_inst_dmem_ram_236__5_), .B(mem_stage_inst_dmem_ram_238__5_), 
        .C(mem_stage_inst_dmem_ram_237__5_), .D(
        mem_stage_inst_dmem_ram_239__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4751) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u751 ( .A(mem_stage_inst_dmem_n4748), 
        .B(mem_stage_inst_dmem_n4749), .C(mem_stage_inst_dmem_n4750), .D(
        mem_stage_inst_dmem_n4751), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4747) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u750 ( .A(mem_stage_inst_dmem_ram_96__5_), .B(mem_stage_inst_dmem_ram_98__5_), .C(mem_stage_inst_dmem_ram_97__5_), .D(
        mem_stage_inst_dmem_ram_99__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4788) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u749 ( .A(
        mem_stage_inst_dmem_ram_100__5_), .B(mem_stage_inst_dmem_ram_102__5_), 
        .C(mem_stage_inst_dmem_ram_101__5_), .D(
        mem_stage_inst_dmem_ram_103__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4790) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u748 ( .A(
        mem_stage_inst_dmem_ram_108__5_), .B(mem_stage_inst_dmem_ram_110__5_), 
        .C(mem_stage_inst_dmem_ram_109__5_), .D(
        mem_stage_inst_dmem_ram_111__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4791) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u747 ( .A(mem_stage_inst_dmem_n4788), 
        .B(mem_stage_inst_dmem_n4789), .C(mem_stage_inst_dmem_n4790), .D(
        mem_stage_inst_dmem_n4791), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4787) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u746 ( .A(mem_stage_inst_dmem_ram_32__5_), .B(mem_stage_inst_dmem_ram_34__5_), .C(mem_stage_inst_dmem_ram_33__5_), .D(
        mem_stage_inst_dmem_ram_35__5_), .S0(mem_stage_inst_dmem_n164), .S1(
        ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4808) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u745 ( .A(mem_stage_inst_dmem_ram_36__5_), .B(mem_stage_inst_dmem_ram_38__5_), .C(mem_stage_inst_dmem_ram_37__5_), .D(
        mem_stage_inst_dmem_ram_39__5_), .S0(mem_stage_inst_dmem_n164), .S1(
        ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4810) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u744 ( .A(mem_stage_inst_dmem_ram_44__5_), .B(mem_stage_inst_dmem_ram_46__5_), .C(mem_stage_inst_dmem_ram_45__5_), .D(
        mem_stage_inst_dmem_ram_47__5_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n4811) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u743 ( .A(mem_stage_inst_dmem_n4808), 
        .B(mem_stage_inst_dmem_n4809), .C(mem_stage_inst_dmem_n4810), .D(
        mem_stage_inst_dmem_n4811), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4807) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u742 ( .A(
        mem_stage_inst_dmem_ram_160__5_), .B(mem_stage_inst_dmem_ram_162__5_), 
        .C(mem_stage_inst_dmem_ram_161__5_), .D(
        mem_stage_inst_dmem_ram_163__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4768) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u741 ( .A(
        mem_stage_inst_dmem_ram_164__5_), .B(mem_stage_inst_dmem_ram_166__5_), 
        .C(mem_stage_inst_dmem_ram_165__5_), .D(
        mem_stage_inst_dmem_ram_167__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4770) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u740 ( .A(
        mem_stage_inst_dmem_ram_172__5_), .B(mem_stage_inst_dmem_ram_174__5_), 
        .C(mem_stage_inst_dmem_ram_173__5_), .D(
        mem_stage_inst_dmem_ram_175__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4771) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u739 ( .A(mem_stage_inst_dmem_n4768), 
        .B(mem_stage_inst_dmem_n4769), .C(mem_stage_inst_dmem_n4770), .D(
        mem_stage_inst_dmem_n4771), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4767) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u738 ( .A(
        mem_stage_inst_dmem_ram_224__4_), .B(mem_stage_inst_dmem_ram_226__4_), 
        .C(mem_stage_inst_dmem_ram_225__4_), .D(
        mem_stage_inst_dmem_ram_227__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4664) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u737 ( .A(
        mem_stage_inst_dmem_ram_228__4_), .B(mem_stage_inst_dmem_ram_230__4_), 
        .C(mem_stage_inst_dmem_ram_229__4_), .D(
        mem_stage_inst_dmem_ram_231__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4666) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u736 ( .A(
        mem_stage_inst_dmem_ram_236__4_), .B(mem_stage_inst_dmem_ram_238__4_), 
        .C(mem_stage_inst_dmem_ram_237__4_), .D(
        mem_stage_inst_dmem_ram_239__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4667) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u735 ( .A(mem_stage_inst_dmem_n4664), 
        .B(mem_stage_inst_dmem_n4665), .C(mem_stage_inst_dmem_n4666), .D(
        mem_stage_inst_dmem_n4667), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4663) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u734 ( .A(mem_stage_inst_dmem_ram_96__4_), .B(mem_stage_inst_dmem_ram_98__4_), .C(mem_stage_inst_dmem_ram_97__4_), .D(
        mem_stage_inst_dmem_ram_99__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4704) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u733 ( .A(
        mem_stage_inst_dmem_ram_100__4_), .B(mem_stage_inst_dmem_ram_102__4_), 
        .C(mem_stage_inst_dmem_ram_101__4_), .D(
        mem_stage_inst_dmem_ram_103__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4706) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u732 ( .A(
        mem_stage_inst_dmem_ram_108__4_), .B(mem_stage_inst_dmem_ram_110__4_), 
        .C(mem_stage_inst_dmem_ram_109__4_), .D(
        mem_stage_inst_dmem_ram_111__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4707) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u731 ( .A(mem_stage_inst_dmem_n4704), 
        .B(mem_stage_inst_dmem_n4705), .C(mem_stage_inst_dmem_n4706), .D(
        mem_stage_inst_dmem_n4707), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4703) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u730 ( .A(mem_stage_inst_dmem_ram_32__4_), .B(mem_stage_inst_dmem_ram_34__4_), .C(mem_stage_inst_dmem_ram_33__4_), .D(
        mem_stage_inst_dmem_ram_35__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4724) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u729 ( .A(mem_stage_inst_dmem_ram_36__4_), .B(mem_stage_inst_dmem_ram_38__4_), .C(mem_stage_inst_dmem_ram_37__4_), .D(
        mem_stage_inst_dmem_ram_39__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4726) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u728 ( .A(mem_stage_inst_dmem_ram_44__4_), .B(mem_stage_inst_dmem_ram_46__4_), .C(mem_stage_inst_dmem_ram_45__4_), .D(
        mem_stage_inst_dmem_ram_47__4_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n4727) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u727 ( .A(mem_stage_inst_dmem_n4724), 
        .B(mem_stage_inst_dmem_n4725), .C(mem_stage_inst_dmem_n4726), .D(
        mem_stage_inst_dmem_n4727), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4723) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u726 ( .A(
        mem_stage_inst_dmem_ram_160__4_), .B(mem_stage_inst_dmem_ram_162__4_), 
        .C(mem_stage_inst_dmem_ram_161__4_), .D(
        mem_stage_inst_dmem_ram_163__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4684) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u725 ( .A(
        mem_stage_inst_dmem_ram_164__4_), .B(mem_stage_inst_dmem_ram_166__4_), 
        .C(mem_stage_inst_dmem_ram_165__4_), .D(
        mem_stage_inst_dmem_ram_167__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4686) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u724 ( .A(
        mem_stage_inst_dmem_ram_172__4_), .B(mem_stage_inst_dmem_ram_174__4_), 
        .C(mem_stage_inst_dmem_ram_173__4_), .D(
        mem_stage_inst_dmem_ram_175__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4687) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u723 ( .A(mem_stage_inst_dmem_n4684), 
        .B(mem_stage_inst_dmem_n4685), .C(mem_stage_inst_dmem_n4686), .D(
        mem_stage_inst_dmem_n4687), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4683) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u722 ( .A(
        mem_stage_inst_dmem_ram_224__3_), .B(mem_stage_inst_dmem_ram_226__3_), 
        .C(mem_stage_inst_dmem_ram_225__3_), .D(
        mem_stage_inst_dmem_ram_227__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n484) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u721 ( .A(
        mem_stage_inst_dmem_ram_228__3_), .B(mem_stage_inst_dmem_ram_230__3_), 
        .C(mem_stage_inst_dmem_ram_229__3_), .D(
        mem_stage_inst_dmem_ram_231__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n486) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u720 ( .A(
        mem_stage_inst_dmem_ram_236__3_), .B(mem_stage_inst_dmem_ram_238__3_), 
        .C(mem_stage_inst_dmem_ram_237__3_), .D(
        mem_stage_inst_dmem_ram_239__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n487) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u719 ( .A(mem_stage_inst_dmem_n484), .B(
        mem_stage_inst_dmem_n485), .C(mem_stage_inst_dmem_n486), .D(
        mem_stage_inst_dmem_n487), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n483) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u718 ( .A(mem_stage_inst_dmem_ram_96__3_), .B(mem_stage_inst_dmem_ram_98__3_), .C(mem_stage_inst_dmem_ram_97__3_), .D(
        mem_stage_inst_dmem_ram_99__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n524) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u717 ( .A(
        mem_stage_inst_dmem_ram_100__3_), .B(mem_stage_inst_dmem_ram_102__3_), 
        .C(mem_stage_inst_dmem_ram_101__3_), .D(
        mem_stage_inst_dmem_ram_103__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n526) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u716 ( .A(
        mem_stage_inst_dmem_ram_108__3_), .B(mem_stage_inst_dmem_ram_110__3_), 
        .C(mem_stage_inst_dmem_ram_109__3_), .D(
        mem_stage_inst_dmem_ram_111__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n527) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u715 ( .A(mem_stage_inst_dmem_n524), .B(
        mem_stage_inst_dmem_n525), .C(mem_stage_inst_dmem_n526), .D(
        mem_stage_inst_dmem_n527), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n523) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u714 ( .A(mem_stage_inst_dmem_ram_32__3_), .B(mem_stage_inst_dmem_ram_34__3_), .C(mem_stage_inst_dmem_ram_33__3_), .D(
        mem_stage_inst_dmem_ram_35__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n544) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u713 ( .A(mem_stage_inst_dmem_ram_36__3_), .B(mem_stage_inst_dmem_ram_38__3_), .C(mem_stage_inst_dmem_ram_37__3_), .D(
        mem_stage_inst_dmem_ram_39__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n546) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u712 ( .A(mem_stage_inst_dmem_ram_44__3_), .B(mem_stage_inst_dmem_ram_46__3_), .C(mem_stage_inst_dmem_ram_45__3_), .D(
        mem_stage_inst_dmem_ram_47__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n547) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u711 ( .A(mem_stage_inst_dmem_n544), .B(
        mem_stage_inst_dmem_n545), .C(mem_stage_inst_dmem_n546), .D(
        mem_stage_inst_dmem_n547), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n543) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u710 ( .A(
        mem_stage_inst_dmem_ram_160__3_), .B(mem_stage_inst_dmem_ram_162__3_), 
        .C(mem_stage_inst_dmem_ram_161__3_), .D(
        mem_stage_inst_dmem_ram_163__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n504) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u709 ( .A(
        mem_stage_inst_dmem_ram_164__3_), .B(mem_stage_inst_dmem_ram_166__3_), 
        .C(mem_stage_inst_dmem_ram_165__3_), .D(
        mem_stage_inst_dmem_ram_167__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n506) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u708 ( .A(
        mem_stage_inst_dmem_ram_172__3_), .B(mem_stage_inst_dmem_ram_174__3_), 
        .C(mem_stage_inst_dmem_ram_173__3_), .D(
        mem_stage_inst_dmem_ram_175__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n507) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u707 ( .A(mem_stage_inst_dmem_n504), .B(
        mem_stage_inst_dmem_n505), .C(mem_stage_inst_dmem_n506), .D(
        mem_stage_inst_dmem_n507), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n503) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u706 ( .A(
        mem_stage_inst_dmem_ram_224__2_), .B(mem_stage_inst_dmem_ram_226__2_), 
        .C(mem_stage_inst_dmem_ram_225__2_), .D(
        mem_stage_inst_dmem_ram_227__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n400) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u705 ( .A(
        mem_stage_inst_dmem_ram_228__2_), .B(mem_stage_inst_dmem_ram_230__2_), 
        .C(mem_stage_inst_dmem_ram_229__2_), .D(
        mem_stage_inst_dmem_ram_231__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n402) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u704 ( .A(
        mem_stage_inst_dmem_ram_236__2_), .B(mem_stage_inst_dmem_ram_238__2_), 
        .C(mem_stage_inst_dmem_ram_237__2_), .D(
        mem_stage_inst_dmem_ram_239__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n403) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u703 ( .A(mem_stage_inst_dmem_n400), .B(
        mem_stage_inst_dmem_n401), .C(mem_stage_inst_dmem_n402), .D(
        mem_stage_inst_dmem_n403), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n399) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u702 ( .A(mem_stage_inst_dmem_ram_96__2_), .B(mem_stage_inst_dmem_ram_98__2_), .C(mem_stage_inst_dmem_ram_97__2_), .D(
        mem_stage_inst_dmem_ram_99__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n440) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u701 ( .A(
        mem_stage_inst_dmem_ram_100__2_), .B(mem_stage_inst_dmem_ram_102__2_), 
        .C(mem_stage_inst_dmem_ram_101__2_), .D(
        mem_stage_inst_dmem_ram_103__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n442) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u700 ( .A(
        mem_stage_inst_dmem_ram_108__2_), .B(mem_stage_inst_dmem_ram_110__2_), 
        .C(mem_stage_inst_dmem_ram_109__2_), .D(
        mem_stage_inst_dmem_ram_111__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n443) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u699 ( .A(mem_stage_inst_dmem_n440), .B(
        mem_stage_inst_dmem_n441), .C(mem_stage_inst_dmem_n442), .D(
        mem_stage_inst_dmem_n443), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n439) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u698 ( .A(mem_stage_inst_dmem_ram_32__2_), .B(mem_stage_inst_dmem_ram_34__2_), .C(mem_stage_inst_dmem_ram_33__2_), .D(
        mem_stage_inst_dmem_ram_35__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n460) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u697 ( .A(mem_stage_inst_dmem_ram_36__2_), .B(mem_stage_inst_dmem_ram_38__2_), .C(mem_stage_inst_dmem_ram_37__2_), .D(
        mem_stage_inst_dmem_ram_39__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n462) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u696 ( .A(mem_stage_inst_dmem_ram_44__2_), .B(mem_stage_inst_dmem_ram_46__2_), .C(mem_stage_inst_dmem_ram_45__2_), .D(
        mem_stage_inst_dmem_ram_47__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n463) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u695 ( .A(mem_stage_inst_dmem_n460), .B(
        mem_stage_inst_dmem_n461), .C(mem_stage_inst_dmem_n462), .D(
        mem_stage_inst_dmem_n463), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n459) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u694 ( .A(
        mem_stage_inst_dmem_ram_160__2_), .B(mem_stage_inst_dmem_ram_162__2_), 
        .C(mem_stage_inst_dmem_ram_161__2_), .D(
        mem_stage_inst_dmem_ram_163__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n420) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u693 ( .A(
        mem_stage_inst_dmem_ram_164__2_), .B(mem_stage_inst_dmem_ram_166__2_), 
        .C(mem_stage_inst_dmem_ram_165__2_), .D(
        mem_stage_inst_dmem_ram_167__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n422) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u692 ( .A(
        mem_stage_inst_dmem_ram_172__2_), .B(mem_stage_inst_dmem_ram_174__2_), 
        .C(mem_stage_inst_dmem_ram_173__2_), .D(
        mem_stage_inst_dmem_ram_175__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n423) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u691 ( .A(mem_stage_inst_dmem_n420), .B(
        mem_stage_inst_dmem_n421), .C(mem_stage_inst_dmem_n422), .D(
        mem_stage_inst_dmem_n423), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n419) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u690 ( .A(
        mem_stage_inst_dmem_ram_224__1_), .B(mem_stage_inst_dmem_ram_226__1_), 
        .C(mem_stage_inst_dmem_ram_225__1_), .D(
        mem_stage_inst_dmem_ram_227__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n316) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u689 ( .A(
        mem_stage_inst_dmem_ram_228__1_), .B(mem_stage_inst_dmem_ram_230__1_), 
        .C(mem_stage_inst_dmem_ram_229__1_), .D(
        mem_stage_inst_dmem_ram_231__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n318) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u688 ( .A(
        mem_stage_inst_dmem_ram_236__1_), .B(mem_stage_inst_dmem_ram_238__1_), 
        .C(mem_stage_inst_dmem_ram_237__1_), .D(
        mem_stage_inst_dmem_ram_239__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n319) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u687 ( .A(mem_stage_inst_dmem_n316), .B(
        mem_stage_inst_dmem_n317), .C(mem_stage_inst_dmem_n318), .D(
        mem_stage_inst_dmem_n319), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n315) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u686 ( .A(mem_stage_inst_dmem_ram_96__1_), .B(mem_stage_inst_dmem_ram_98__1_), .C(mem_stage_inst_dmem_ram_97__1_), .D(
        mem_stage_inst_dmem_ram_99__1_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n356) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u685 ( .A(
        mem_stage_inst_dmem_ram_100__1_), .B(mem_stage_inst_dmem_ram_102__1_), 
        .C(mem_stage_inst_dmem_ram_101__1_), .D(
        mem_stage_inst_dmem_ram_103__1_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n358) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u684 ( .A(
        mem_stage_inst_dmem_ram_108__1_), .B(mem_stage_inst_dmem_ram_110__1_), 
        .C(mem_stage_inst_dmem_ram_109__1_), .D(
        mem_stage_inst_dmem_ram_111__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n359) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u683 ( .A(mem_stage_inst_dmem_n356), .B(
        mem_stage_inst_dmem_n357), .C(mem_stage_inst_dmem_n358), .D(
        mem_stage_inst_dmem_n359), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n355) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u682 ( .A(mem_stage_inst_dmem_ram_32__1_), .B(mem_stage_inst_dmem_ram_34__1_), .C(mem_stage_inst_dmem_ram_33__1_), .D(
        mem_stage_inst_dmem_ram_35__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n376) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u681 ( .A(mem_stage_inst_dmem_ram_36__1_), .B(mem_stage_inst_dmem_ram_38__1_), .C(mem_stage_inst_dmem_ram_37__1_), .D(
        mem_stage_inst_dmem_ram_39__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n378) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u680 ( .A(mem_stage_inst_dmem_ram_44__1_), .B(mem_stage_inst_dmem_ram_46__1_), .C(mem_stage_inst_dmem_ram_45__1_), .D(
        mem_stage_inst_dmem_ram_47__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n379) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u679 ( .A(mem_stage_inst_dmem_n376), .B(
        mem_stage_inst_dmem_n377), .C(mem_stage_inst_dmem_n378), .D(
        mem_stage_inst_dmem_n379), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n375) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u678 ( .A(
        mem_stage_inst_dmem_ram_160__1_), .B(mem_stage_inst_dmem_ram_162__1_), 
        .C(mem_stage_inst_dmem_ram_161__1_), .D(
        mem_stage_inst_dmem_ram_163__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n336) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u677 ( .A(
        mem_stage_inst_dmem_ram_164__1_), .B(mem_stage_inst_dmem_ram_166__1_), 
        .C(mem_stage_inst_dmem_ram_165__1_), .D(
        mem_stage_inst_dmem_ram_167__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n338) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u676 ( .A(
        mem_stage_inst_dmem_ram_172__1_), .B(mem_stage_inst_dmem_ram_174__1_), 
        .C(mem_stage_inst_dmem_ram_173__1_), .D(
        mem_stage_inst_dmem_ram_175__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n339) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u675 ( .A(mem_stage_inst_dmem_n336), .B(
        mem_stage_inst_dmem_n337), .C(mem_stage_inst_dmem_n338), .D(
        mem_stage_inst_dmem_n339), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n335) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u674 ( .A(
        mem_stage_inst_dmem_ram_224__0_), .B(mem_stage_inst_dmem_ram_226__0_), 
        .C(mem_stage_inst_dmem_ram_225__0_), .D(
        mem_stage_inst_dmem_ram_227__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n232) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u673 ( .A(
        mem_stage_inst_dmem_ram_228__0_), .B(mem_stage_inst_dmem_ram_230__0_), 
        .C(mem_stage_inst_dmem_ram_229__0_), .D(
        mem_stage_inst_dmem_ram_231__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n234) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u672 ( .A(
        mem_stage_inst_dmem_ram_236__0_), .B(mem_stage_inst_dmem_ram_238__0_), 
        .C(mem_stage_inst_dmem_ram_237__0_), .D(
        mem_stage_inst_dmem_ram_239__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n235) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u671 ( .A(mem_stage_inst_dmem_n232), .B(
        mem_stage_inst_dmem_n233), .C(mem_stage_inst_dmem_n234), .D(
        mem_stage_inst_dmem_n235), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n231) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u670 ( .A(mem_stage_inst_dmem_ram_96__0_), .B(mem_stage_inst_dmem_ram_98__0_), .C(mem_stage_inst_dmem_ram_97__0_), .D(
        mem_stage_inst_dmem_ram_99__0_), .S0(mem_stage_inst_dmem_n138), .S1(
        mem_stage_inst_dmem_n40), .Y(mem_stage_inst_dmem_n272) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u669 ( .A(
        mem_stage_inst_dmem_ram_100__0_), .B(mem_stage_inst_dmem_ram_102__0_), 
        .C(mem_stage_inst_dmem_ram_101__0_), .D(
        mem_stage_inst_dmem_ram_103__0_), .S0(mem_stage_inst_dmem_n138), .S1(
        mem_stage_inst_dmem_n40), .Y(mem_stage_inst_dmem_n274) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u668 ( .A(
        mem_stage_inst_dmem_ram_108__0_), .B(mem_stage_inst_dmem_ram_110__0_), 
        .C(mem_stage_inst_dmem_ram_109__0_), .D(
        mem_stage_inst_dmem_ram_111__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n275) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u667 ( .A(mem_stage_inst_dmem_n272), .B(
        mem_stage_inst_dmem_n273), .C(mem_stage_inst_dmem_n274), .D(
        mem_stage_inst_dmem_n275), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n271) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u666 ( .A(mem_stage_inst_dmem_ram_32__0_), .B(mem_stage_inst_dmem_ram_34__0_), .C(mem_stage_inst_dmem_ram_33__0_), .D(
        mem_stage_inst_dmem_ram_35__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n292) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u665 ( .A(mem_stage_inst_dmem_ram_36__0_), .B(mem_stage_inst_dmem_ram_38__0_), .C(mem_stage_inst_dmem_ram_37__0_), .D(
        mem_stage_inst_dmem_ram_39__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n294) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u664 ( .A(mem_stage_inst_dmem_ram_44__0_), .B(mem_stage_inst_dmem_ram_46__0_), .C(mem_stage_inst_dmem_ram_45__0_), .D(
        mem_stage_inst_dmem_ram_47__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n295) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u663 ( .A(mem_stage_inst_dmem_n292), .B(
        mem_stage_inst_dmem_n293), .C(mem_stage_inst_dmem_n294), .D(
        mem_stage_inst_dmem_n295), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n291) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u662 ( .A(
        mem_stage_inst_dmem_ram_160__0_), .B(mem_stage_inst_dmem_ram_162__0_), 
        .C(mem_stage_inst_dmem_ram_161__0_), .D(
        mem_stage_inst_dmem_ram_163__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n252) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u661 ( .A(
        mem_stage_inst_dmem_ram_164__0_), .B(mem_stage_inst_dmem_ram_166__0_), 
        .C(mem_stage_inst_dmem_ram_165__0_), .D(
        mem_stage_inst_dmem_ram_167__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n254) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u660 ( .A(
        mem_stage_inst_dmem_ram_172__0_), .B(mem_stage_inst_dmem_ram_174__0_), 
        .C(mem_stage_inst_dmem_ram_173__0_), .D(
        mem_stage_inst_dmem_ram_175__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n255) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u659 ( .A(mem_stage_inst_dmem_n252), .B(
        mem_stage_inst_dmem_n253), .C(mem_stage_inst_dmem_n254), .D(
        mem_stage_inst_dmem_n255), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n251) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u658 ( .A(
        mem_stage_inst_dmem_ram_248__15_), .B(mem_stage_inst_dmem_ram_250__15_), .C(mem_stage_inst_dmem_ram_249__15_), .D(mem_stage_inst_dmem_ram_251__15_), 
        .S0(mem_stage_inst_dmem_n139), .S1(mem_stage_inst_dmem_n29), .Y(
        mem_stage_inst_dmem_n5584) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u657 ( .A(
        mem_stage_inst_dmem_ram_216__15_), .B(mem_stage_inst_dmem_ram_218__15_), .C(mem_stage_inst_dmem_ram_217__15_), .D(mem_stage_inst_dmem_ram_219__15_), 
        .S0(mem_stage_inst_dmem_n150), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5594) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u656 ( .A(
        mem_stage_inst_dmem_ram_200__15_), .B(mem_stage_inst_dmem_ram_202__15_), .C(mem_stage_inst_dmem_ram_201__15_), .D(mem_stage_inst_dmem_ram_203__15_), 
        .S0(mem_stage_inst_dmem_n148), .S1(mem_stage_inst_dmem_n61), .Y(
        mem_stage_inst_dmem_n5599) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u655 ( .A(
        mem_stage_inst_dmem_ram_232__15_), .B(mem_stage_inst_dmem_ram_234__15_), .C(mem_stage_inst_dmem_ram_233__15_), .D(mem_stage_inst_dmem_ram_235__15_), 
        .S0(mem_stage_inst_dmem_n149), .S1(mem_stage_inst_dmem_n62), .Y(
        mem_stage_inst_dmem_n5589) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u654 ( .A(
        mem_stage_inst_dmem_ram_120__15_), .B(mem_stage_inst_dmem_ram_122__15_), .C(mem_stage_inst_dmem_ram_121__15_), .D(mem_stage_inst_dmem_ram_123__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n33), .Y(
        mem_stage_inst_dmem_n5624) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u653 ( .A(
        mem_stage_inst_dmem_ram_88__15_), .B(mem_stage_inst_dmem_ram_90__15_), 
        .C(mem_stage_inst_dmem_ram_89__15_), .D(
        mem_stage_inst_dmem_ram_91__15_), .S0(ex_pipeline_reg_out[23]), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n5634) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u652 ( .A(
        mem_stage_inst_dmem_ram_72__15_), .B(mem_stage_inst_dmem_ram_74__15_), 
        .C(mem_stage_inst_dmem_ram_73__15_), .D(
        mem_stage_inst_dmem_ram_75__15_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n50), .Y(mem_stage_inst_dmem_n5639) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u651 ( .A(
        mem_stage_inst_dmem_ram_104__15_), .B(mem_stage_inst_dmem_ram_106__15_), .C(mem_stage_inst_dmem_ram_105__15_), .D(mem_stage_inst_dmem_ram_107__15_), 
        .S0(ex_pipeline_reg_out[23]), .S1(mem_stage_inst_dmem_n38), .Y(
        mem_stage_inst_dmem_n5629) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u650 ( .A(
        mem_stage_inst_dmem_ram_56__15_), .B(mem_stage_inst_dmem_ram_58__15_), 
        .C(mem_stage_inst_dmem_ram_57__15_), .D(
        mem_stage_inst_dmem_ram_59__15_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5644) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u649 ( .A(
        mem_stage_inst_dmem_ram_24__15_), .B(mem_stage_inst_dmem_ram_26__15_), 
        .C(mem_stage_inst_dmem_ram_25__15_), .D(
        mem_stage_inst_dmem_ram_27__15_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n5654) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u648 ( .A(mem_stage_inst_dmem_ram_8__15_), .B(mem_stage_inst_dmem_ram_10__15_), .C(mem_stage_inst_dmem_ram_9__15_), .D(
        mem_stage_inst_dmem_ram_11__15_), .S0(mem_stage_inst_dmem_n116), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n5659) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u647 ( .A(
        mem_stage_inst_dmem_ram_40__15_), .B(mem_stage_inst_dmem_ram_42__15_), 
        .C(mem_stage_inst_dmem_ram_41__15_), .D(
        mem_stage_inst_dmem_ram_43__15_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n5649) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u646 ( .A(
        mem_stage_inst_dmem_ram_184__15_), .B(mem_stage_inst_dmem_ram_186__15_), .C(mem_stage_inst_dmem_ram_185__15_), .D(mem_stage_inst_dmem_ram_187__15_), 
        .S0(mem_stage_inst_dmem_n159), .S1(mem_stage_inst_dmem_n9), .Y(
        mem_stage_inst_dmem_n5604) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u645 ( .A(
        mem_stage_inst_dmem_ram_152__15_), .B(mem_stage_inst_dmem_ram_154__15_), .C(mem_stage_inst_dmem_ram_153__15_), .D(mem_stage_inst_dmem_ram_155__15_), 
        .S0(mem_stage_inst_dmem_n157), .S1(mem_stage_inst_dmem_n10), .Y(
        mem_stage_inst_dmem_n5614) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u644 ( .A(
        mem_stage_inst_dmem_ram_136__15_), .B(mem_stage_inst_dmem_ram_138__15_), .C(mem_stage_inst_dmem_ram_137__15_), .D(mem_stage_inst_dmem_ram_139__15_), 
        .S0(mem_stage_inst_dmem_n158), .S1(mem_stage_inst_dmem_n11), .Y(
        mem_stage_inst_dmem_n5619) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u643 ( .A(
        mem_stage_inst_dmem_ram_168__15_), .B(mem_stage_inst_dmem_ram_170__15_), .C(mem_stage_inst_dmem_ram_169__15_), .D(mem_stage_inst_dmem_ram_171__15_), 
        .S0(mem_stage_inst_dmem_n160), .S1(mem_stage_inst_dmem_n13), .Y(
        mem_stage_inst_dmem_n5609) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u642 ( .A(
        mem_stage_inst_dmem_ram_248__14_), .B(mem_stage_inst_dmem_ram_250__14_), .C(mem_stage_inst_dmem_ram_249__14_), .D(mem_stage_inst_dmem_ram_251__14_), 
        .S0(mem_stage_inst_dmem_n156), .S1(mem_stage_inst_dmem_n64), .Y(
        mem_stage_inst_dmem_n5500) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u641 ( .A(
        mem_stage_inst_dmem_ram_216__14_), .B(mem_stage_inst_dmem_ram_218__14_), .C(mem_stage_inst_dmem_ram_217__14_), .D(mem_stage_inst_dmem_ram_219__14_), 
        .S0(mem_stage_inst_dmem_n135), .S1(mem_stage_inst_dmem_n57), .Y(
        mem_stage_inst_dmem_n5510) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u640 ( .A(
        mem_stage_inst_dmem_ram_200__14_), .B(mem_stage_inst_dmem_ram_202__14_), .C(mem_stage_inst_dmem_ram_201__14_), .D(mem_stage_inst_dmem_ram_203__14_), 
        .S0(mem_stage_inst_dmem_n133), .S1(mem_stage_inst_dmem_n50), .Y(
        mem_stage_inst_dmem_n5515) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u639 ( .A(
        mem_stage_inst_dmem_ram_232__14_), .B(mem_stage_inst_dmem_ram_234__14_), .C(mem_stage_inst_dmem_ram_233__14_), .D(mem_stage_inst_dmem_ram_235__14_), 
        .S0(mem_stage_inst_dmem_n134), .S1(mem_stage_inst_dmem_n51), .Y(
        mem_stage_inst_dmem_n5505) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u638 ( .A(
        mem_stage_inst_dmem_ram_120__14_), .B(mem_stage_inst_dmem_ram_122__14_), .C(mem_stage_inst_dmem_ram_121__14_), .D(mem_stage_inst_dmem_ram_123__14_), 
        .S0(mem_stage_inst_dmem_n153), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5540) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u637 ( .A(
        mem_stage_inst_dmem_ram_88__14_), .B(mem_stage_inst_dmem_ram_90__14_), 
        .C(mem_stage_inst_dmem_ram_89__14_), .D(
        mem_stage_inst_dmem_ram_91__14_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5550) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u636 ( .A(
        mem_stage_inst_dmem_ram_72__14_), .B(mem_stage_inst_dmem_ram_74__14_), 
        .C(mem_stage_inst_dmem_ram_73__14_), .D(
        mem_stage_inst_dmem_ram_75__14_), .S0(mem_stage_inst_dmem_n118), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5555) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u635 ( .A(
        mem_stage_inst_dmem_ram_104__14_), .B(mem_stage_inst_dmem_ram_106__14_), .C(mem_stage_inst_dmem_ram_105__14_), .D(mem_stage_inst_dmem_ram_107__14_), 
        .S0(mem_stage_inst_dmem_n155), .S1(mem_stage_inst_dmem_n20), .Y(
        mem_stage_inst_dmem_n5545) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u634 ( .A(
        mem_stage_inst_dmem_ram_56__14_), .B(mem_stage_inst_dmem_ram_58__14_), 
        .C(mem_stage_inst_dmem_ram_57__14_), .D(
        mem_stage_inst_dmem_ram_59__14_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5560) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u633 ( .A(
        mem_stage_inst_dmem_ram_24__14_), .B(mem_stage_inst_dmem_ram_26__14_), 
        .C(mem_stage_inst_dmem_ram_25__14_), .D(
        mem_stage_inst_dmem_ram_27__14_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n5570) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u632 ( .A(mem_stage_inst_dmem_ram_8__14_), .B(mem_stage_inst_dmem_ram_10__14_), .C(mem_stage_inst_dmem_ram_9__14_), .D(
        mem_stage_inst_dmem_ram_11__14_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n5575) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u631 ( .A(
        mem_stage_inst_dmem_ram_40__14_), .B(mem_stage_inst_dmem_ram_42__14_), 
        .C(mem_stage_inst_dmem_ram_41__14_), .D(
        mem_stage_inst_dmem_ram_43__14_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5565) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u630 ( .A(
        mem_stage_inst_dmem_ram_184__14_), .B(mem_stage_inst_dmem_ram_186__14_), .C(mem_stage_inst_dmem_ram_185__14_), .D(mem_stage_inst_dmem_ram_187__14_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5520) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u629 ( .A(
        mem_stage_inst_dmem_ram_152__14_), .B(mem_stage_inst_dmem_ram_154__14_), .C(mem_stage_inst_dmem_ram_153__14_), .D(mem_stage_inst_dmem_ram_155__14_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5530) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u628 ( .A(
        mem_stage_inst_dmem_ram_136__14_), .B(mem_stage_inst_dmem_ram_138__14_), .C(mem_stage_inst_dmem_ram_137__14_), .D(mem_stage_inst_dmem_ram_139__14_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5535) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u627 ( .A(
        mem_stage_inst_dmem_ram_168__14_), .B(mem_stage_inst_dmem_ram_170__14_), .C(mem_stage_inst_dmem_ram_169__14_), .D(mem_stage_inst_dmem_ram_171__14_), 
        .S0(mem_stage_inst_dmem_n124), .S1(mem_stage_inst_dmem_n19), .Y(
        mem_stage_inst_dmem_n5525) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u626 ( .A(
        mem_stage_inst_dmem_ram_248__13_), .B(mem_stage_inst_dmem_ram_250__13_), .C(mem_stage_inst_dmem_ram_249__13_), .D(mem_stage_inst_dmem_ram_251__13_), 
        .S0(mem_stage_inst_dmem_n142), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5416) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u625 ( .A(
        mem_stage_inst_dmem_ram_216__13_), .B(mem_stage_inst_dmem_ram_218__13_), .C(mem_stage_inst_dmem_ram_217__13_), .D(mem_stage_inst_dmem_ram_219__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5426) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u624 ( .A(
        mem_stage_inst_dmem_ram_200__13_), .B(mem_stage_inst_dmem_ram_202__13_), .C(mem_stage_inst_dmem_ram_201__13_), .D(mem_stage_inst_dmem_ram_203__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5431) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u623 ( .A(
        mem_stage_inst_dmem_ram_232__13_), .B(mem_stage_inst_dmem_ram_234__13_), .C(mem_stage_inst_dmem_ram_233__13_), .D(mem_stage_inst_dmem_ram_235__13_), 
        .S0(mem_stage_inst_dmem_n143), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5421) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u622 ( .A(
        mem_stage_inst_dmem_ram_120__13_), .B(mem_stage_inst_dmem_ram_122__13_), .C(mem_stage_inst_dmem_ram_121__13_), .D(mem_stage_inst_dmem_ram_123__13_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n53), .Y(
        mem_stage_inst_dmem_n5456) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u621 ( .A(
        mem_stage_inst_dmem_ram_88__13_), .B(mem_stage_inst_dmem_ram_90__13_), 
        .C(mem_stage_inst_dmem_ram_89__13_), .D(
        mem_stage_inst_dmem_ram_91__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n5466) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u620 ( .A(
        mem_stage_inst_dmem_ram_72__13_), .B(mem_stage_inst_dmem_ram_74__13_), 
        .C(mem_stage_inst_dmem_ram_73__13_), .D(
        mem_stage_inst_dmem_ram_75__13_), .S0(mem_stage_inst_dmem_n123), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n5471) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u619 ( .A(
        mem_stage_inst_dmem_ram_104__13_), .B(mem_stage_inst_dmem_ram_106__13_), .C(mem_stage_inst_dmem_ram_105__13_), .D(mem_stage_inst_dmem_ram_107__13_), 
        .S0(mem_stage_inst_dmem_n123), .S1(mem_stage_inst_dmem_n56), .Y(
        mem_stage_inst_dmem_n5461) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u618 ( .A(
        mem_stage_inst_dmem_ram_56__13_), .B(mem_stage_inst_dmem_ram_58__13_), 
        .C(mem_stage_inst_dmem_ram_57__13_), .D(
        mem_stage_inst_dmem_ram_59__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5476) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u617 ( .A(
        mem_stage_inst_dmem_ram_24__13_), .B(mem_stage_inst_dmem_ram_26__13_), 
        .C(mem_stage_inst_dmem_ram_25__13_), .D(
        mem_stage_inst_dmem_ram_27__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5486) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u616 ( .A(mem_stage_inst_dmem_ram_8__13_), .B(mem_stage_inst_dmem_ram_10__13_), .C(mem_stage_inst_dmem_ram_9__13_), .D(
        mem_stage_inst_dmem_ram_11__13_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n5491) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u615 ( .A(
        mem_stage_inst_dmem_ram_40__13_), .B(mem_stage_inst_dmem_ram_42__13_), 
        .C(mem_stage_inst_dmem_ram_41__13_), .D(
        mem_stage_inst_dmem_ram_43__13_), .S0(mem_stage_inst_dmem_n124), .S1(
        mem_stage_inst_dmem_n26), .Y(mem_stage_inst_dmem_n5481) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u614 ( .A(
        mem_stage_inst_dmem_ram_184__13_), .B(mem_stage_inst_dmem_ram_186__13_), .C(mem_stage_inst_dmem_ram_185__13_), .D(mem_stage_inst_dmem_ram_187__13_), 
        .S0(mem_stage_inst_dmem_n121), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5436) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u613 ( .A(
        mem_stage_inst_dmem_ram_152__13_), .B(mem_stage_inst_dmem_ram_154__13_), .C(mem_stage_inst_dmem_ram_153__13_), .D(mem_stage_inst_dmem_ram_155__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5446) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u612 ( .A(
        mem_stage_inst_dmem_ram_136__13_), .B(mem_stage_inst_dmem_ram_138__13_), .C(mem_stage_inst_dmem_ram_137__13_), .D(mem_stage_inst_dmem_ram_139__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5451) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u611 ( .A(
        mem_stage_inst_dmem_ram_168__13_), .B(mem_stage_inst_dmem_ram_170__13_), .C(mem_stage_inst_dmem_ram_169__13_), .D(mem_stage_inst_dmem_ram_171__13_), 
        .S0(mem_stage_inst_dmem_n122), .S1(mem_stage_inst_dmem_n25), .Y(
        mem_stage_inst_dmem_n5441) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u610 ( .A(
        mem_stage_inst_dmem_ram_248__12_), .B(mem_stage_inst_dmem_ram_250__12_), .C(mem_stage_inst_dmem_ram_249__12_), .D(mem_stage_inst_dmem_ram_251__12_), 
        .S0(mem_stage_inst_dmem_n116), .S1(mem_stage_inst_dmem_n42), .Y(
        mem_stage_inst_dmem_n5332) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u609 ( .A(
        mem_stage_inst_dmem_ram_216__12_), .B(mem_stage_inst_dmem_ram_218__12_), .C(mem_stage_inst_dmem_ram_217__12_), .D(mem_stage_inst_dmem_ram_219__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5342) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u608 ( .A(
        mem_stage_inst_dmem_ram_200__12_), .B(mem_stage_inst_dmem_ram_202__12_), .C(mem_stage_inst_dmem_ram_201__12_), .D(mem_stage_inst_dmem_ram_203__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5347) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u607 ( .A(
        mem_stage_inst_dmem_ram_232__12_), .B(mem_stage_inst_dmem_ram_234__12_), .C(mem_stage_inst_dmem_ram_233__12_), .D(mem_stage_inst_dmem_ram_235__12_), 
        .S0(mem_stage_inst_dmem_n125), .S1(mem_stage_inst_dmem_n43), .Y(
        mem_stage_inst_dmem_n5337) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u606 ( .A(
        mem_stage_inst_dmem_ram_120__12_), .B(mem_stage_inst_dmem_ram_122__12_), .C(mem_stage_inst_dmem_ram_121__12_), .D(mem_stage_inst_dmem_ram_123__12_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5372) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u605 ( .A(
        mem_stage_inst_dmem_ram_88__12_), .B(mem_stage_inst_dmem_ram_90__12_), 
        .C(mem_stage_inst_dmem_ram_89__12_), .D(
        mem_stage_inst_dmem_ram_91__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5382) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u604 ( .A(
        mem_stage_inst_dmem_ram_72__12_), .B(mem_stage_inst_dmem_ram_74__12_), 
        .C(mem_stage_inst_dmem_ram_73__12_), .D(
        mem_stage_inst_dmem_ram_75__12_), .S0(mem_stage_inst_dmem_n119), .S1(
        mem_stage_inst_dmem_n24), .Y(mem_stage_inst_dmem_n5387) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u603 ( .A(
        mem_stage_inst_dmem_ram_104__12_), .B(mem_stage_inst_dmem_ram_106__12_), .C(mem_stage_inst_dmem_ram_105__12_), .D(mem_stage_inst_dmem_ram_107__12_), 
        .S0(mem_stage_inst_dmem_n119), .S1(mem_stage_inst_dmem_n24), .Y(
        mem_stage_inst_dmem_n5377) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u602 ( .A(
        mem_stage_inst_dmem_ram_56__12_), .B(mem_stage_inst_dmem_ram_58__12_), 
        .C(mem_stage_inst_dmem_ram_57__12_), .D(
        mem_stage_inst_dmem_ram_59__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n5392) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u601 ( .A(
        mem_stage_inst_dmem_ram_24__12_), .B(mem_stage_inst_dmem_ram_26__12_), 
        .C(mem_stage_inst_dmem_ram_25__12_), .D(
        mem_stage_inst_dmem_ram_27__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n20), .Y(mem_stage_inst_dmem_n5402) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u600 ( .A(mem_stage_inst_dmem_ram_8__12_), .B(mem_stage_inst_dmem_ram_10__12_), .C(mem_stage_inst_dmem_ram_9__12_), .D(
        mem_stage_inst_dmem_ram_11__12_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5407) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u599 ( .A(
        mem_stage_inst_dmem_ram_40__12_), .B(mem_stage_inst_dmem_ram_42__12_), 
        .C(mem_stage_inst_dmem_ram_41__12_), .D(
        mem_stage_inst_dmem_ram_43__12_), .S0(mem_stage_inst_dmem_n120), .S1(
        mem_stage_inst_dmem_n21), .Y(mem_stage_inst_dmem_n5397) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u598 ( .A(
        mem_stage_inst_dmem_ram_184__12_), .B(mem_stage_inst_dmem_ram_186__12_), .C(mem_stage_inst_dmem_ram_185__12_), .D(mem_stage_inst_dmem_ram_187__12_), 
        .S0(mem_stage_inst_dmem_n117), .S1(mem_stage_inst_dmem_n22), .Y(
        mem_stage_inst_dmem_n5352) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u597 ( .A(
        mem_stage_inst_dmem_ram_152__12_), .B(mem_stage_inst_dmem_ram_154__12_), .C(mem_stage_inst_dmem_ram_153__12_), .D(mem_stage_inst_dmem_ram_155__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5362) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u596 ( .A(
        mem_stage_inst_dmem_ram_136__12_), .B(mem_stage_inst_dmem_ram_138__12_), .C(mem_stage_inst_dmem_ram_137__12_), .D(mem_stage_inst_dmem_ram_139__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5367) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u595 ( .A(
        mem_stage_inst_dmem_ram_168__12_), .B(mem_stage_inst_dmem_ram_170__12_), .C(mem_stage_inst_dmem_ram_169__12_), .D(mem_stage_inst_dmem_ram_171__12_), 
        .S0(mem_stage_inst_dmem_n118), .S1(mem_stage_inst_dmem_n23), .Y(
        mem_stage_inst_dmem_n5357) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u594 ( .A(
        mem_stage_inst_dmem_ram_248__11_), .B(mem_stage_inst_dmem_ram_250__11_), .C(mem_stage_inst_dmem_ram_249__11_), .D(mem_stage_inst_dmem_ram_251__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5248) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u593 ( .A(
        mem_stage_inst_dmem_ram_216__11_), .B(mem_stage_inst_dmem_ram_218__11_), .C(mem_stage_inst_dmem_ram_217__11_), .D(mem_stage_inst_dmem_ram_219__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5258) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u592 ( .A(
        mem_stage_inst_dmem_ram_200__11_), .B(mem_stage_inst_dmem_ram_202__11_), .C(mem_stage_inst_dmem_ram_201__11_), .D(mem_stage_inst_dmem_ram_203__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5263) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u591 ( .A(
        mem_stage_inst_dmem_ram_232__11_), .B(mem_stage_inst_dmem_ram_234__11_), .C(mem_stage_inst_dmem_ram_233__11_), .D(mem_stage_inst_dmem_ram_235__11_), 
        .S0(mem_stage_inst_dmem_n104), .S1(mem_stage_inst_dmem_n6), .Y(
        mem_stage_inst_dmem_n5253) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u590 ( .A(
        mem_stage_inst_dmem_ram_120__11_), .B(mem_stage_inst_dmem_ram_122__11_), .C(mem_stage_inst_dmem_ram_121__11_), .D(mem_stage_inst_dmem_ram_123__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5288) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u589 ( .A(
        mem_stage_inst_dmem_ram_88__11_), .B(mem_stage_inst_dmem_ram_90__11_), 
        .C(mem_stage_inst_dmem_ram_89__11_), .D(
        mem_stage_inst_dmem_ram_91__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5298) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u588 ( .A(
        mem_stage_inst_dmem_ram_72__11_), .B(mem_stage_inst_dmem_ram_74__11_), 
        .C(mem_stage_inst_dmem_ram_73__11_), .D(
        mem_stage_inst_dmem_ram_75__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5303) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u587 ( .A(
        mem_stage_inst_dmem_ram_104__11_), .B(mem_stage_inst_dmem_ram_106__11_), .C(mem_stage_inst_dmem_ram_105__11_), .D(mem_stage_inst_dmem_ram_107__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5293) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u586 ( .A(
        mem_stage_inst_dmem_ram_56__11_), .B(mem_stage_inst_dmem_ram_58__11_), 
        .C(mem_stage_inst_dmem_ram_57__11_), .D(
        mem_stage_inst_dmem_ram_59__11_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n9), .Y(mem_stage_inst_dmem_n5308) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u585 ( .A(
        mem_stage_inst_dmem_ram_24__11_), .B(mem_stage_inst_dmem_ram_26__11_), 
        .C(mem_stage_inst_dmem_ram_25__11_), .D(
        mem_stage_inst_dmem_ram_27__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5318) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u584 ( .A(mem_stage_inst_dmem_ram_8__11_), .B(mem_stage_inst_dmem_ram_10__11_), .C(mem_stage_inst_dmem_ram_9__11_), .D(
        mem_stage_inst_dmem_ram_11__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5323) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u583 ( .A(
        mem_stage_inst_dmem_ram_40__11_), .B(mem_stage_inst_dmem_ram_42__11_), 
        .C(mem_stage_inst_dmem_ram_41__11_), .D(
        mem_stage_inst_dmem_ram_43__11_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n10), .Y(mem_stage_inst_dmem_n5313) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u582 ( .A(
        mem_stage_inst_dmem_ram_184__11_), .B(mem_stage_inst_dmem_ram_186__11_), .C(mem_stage_inst_dmem_ram_185__11_), .D(mem_stage_inst_dmem_ram_187__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5268) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u581 ( .A(
        mem_stage_inst_dmem_ram_152__11_), .B(mem_stage_inst_dmem_ram_154__11_), .C(mem_stage_inst_dmem_ram_153__11_), .D(mem_stage_inst_dmem_ram_155__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5278) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u580 ( .A(
        mem_stage_inst_dmem_ram_136__11_), .B(mem_stage_inst_dmem_ram_138__11_), .C(mem_stage_inst_dmem_ram_137__11_), .D(mem_stage_inst_dmem_ram_139__11_), 
        .S0(mem_stage_inst_dmem_n106), .S1(mem_stage_inst_dmem_n8), .Y(
        mem_stage_inst_dmem_n5283) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u579 ( .A(
        mem_stage_inst_dmem_ram_168__11_), .B(mem_stage_inst_dmem_ram_170__11_), .C(mem_stage_inst_dmem_ram_169__11_), .D(mem_stage_inst_dmem_ram_171__11_), 
        .S0(mem_stage_inst_dmem_n105), .S1(mem_stage_inst_dmem_n7), .Y(
        mem_stage_inst_dmem_n5273) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u578 ( .A(
        mem_stage_inst_dmem_ram_248__10_), .B(mem_stage_inst_dmem_ram_250__10_), .C(mem_stage_inst_dmem_ram_249__10_), .D(mem_stage_inst_dmem_ram_251__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5164) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u577 ( .A(
        mem_stage_inst_dmem_ram_216__10_), .B(mem_stage_inst_dmem_ram_218__10_), .C(mem_stage_inst_dmem_ram_217__10_), .D(mem_stage_inst_dmem_ram_219__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5174) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u576 ( .A(
        mem_stage_inst_dmem_ram_200__10_), .B(mem_stage_inst_dmem_ram_202__10_), .C(mem_stage_inst_dmem_ram_201__10_), .D(mem_stage_inst_dmem_ram_203__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5179) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u575 ( .A(
        mem_stage_inst_dmem_ram_232__10_), .B(mem_stage_inst_dmem_ram_234__10_), .C(mem_stage_inst_dmem_ram_233__10_), .D(mem_stage_inst_dmem_ram_235__10_), 
        .S0(mem_stage_inst_dmem_n99), .S1(mem_stage_inst_dmem_n1), .Y(
        mem_stage_inst_dmem_n5169) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u574 ( .A(
        mem_stage_inst_dmem_ram_120__10_), .B(mem_stage_inst_dmem_ram_122__10_), .C(mem_stage_inst_dmem_ram_121__10_), .D(mem_stage_inst_dmem_ram_123__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5204) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u573 ( .A(
        mem_stage_inst_dmem_ram_88__10_), .B(mem_stage_inst_dmem_ram_90__10_), 
        .C(mem_stage_inst_dmem_ram_89__10_), .D(
        mem_stage_inst_dmem_ram_91__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5214) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u572 ( .A(
        mem_stage_inst_dmem_ram_72__10_), .B(mem_stage_inst_dmem_ram_74__10_), 
        .C(mem_stage_inst_dmem_ram_73__10_), .D(
        mem_stage_inst_dmem_ram_75__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5219) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u571 ( .A(
        mem_stage_inst_dmem_ram_104__10_), .B(mem_stage_inst_dmem_ram_106__10_), .C(mem_stage_inst_dmem_ram_105__10_), .D(mem_stage_inst_dmem_ram_107__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5209) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u570 ( .A(
        mem_stage_inst_dmem_ram_56__10_), .B(mem_stage_inst_dmem_ram_58__10_), 
        .C(mem_stage_inst_dmem_ram_57__10_), .D(
        mem_stage_inst_dmem_ram_59__10_), .S0(mem_stage_inst_dmem_n102), .S1(
        mem_stage_inst_dmem_n4), .Y(mem_stage_inst_dmem_n5224) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u569 ( .A(
        mem_stage_inst_dmem_ram_24__10_), .B(mem_stage_inst_dmem_ram_26__10_), 
        .C(mem_stage_inst_dmem_ram_25__10_), .D(
        mem_stage_inst_dmem_ram_27__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5234) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u568 ( .A(mem_stage_inst_dmem_ram_8__10_), .B(mem_stage_inst_dmem_ram_10__10_), .C(mem_stage_inst_dmem_ram_9__10_), .D(
        mem_stage_inst_dmem_ram_11__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5239) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u567 ( .A(
        mem_stage_inst_dmem_ram_40__10_), .B(mem_stage_inst_dmem_ram_42__10_), 
        .C(mem_stage_inst_dmem_ram_41__10_), .D(
        mem_stage_inst_dmem_ram_43__10_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n5), .Y(mem_stage_inst_dmem_n5229) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u566 ( .A(
        mem_stage_inst_dmem_ram_184__10_), .B(mem_stage_inst_dmem_ram_186__10_), .C(mem_stage_inst_dmem_ram_185__10_), .D(mem_stage_inst_dmem_ram_187__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5184) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u565 ( .A(
        mem_stage_inst_dmem_ram_152__10_), .B(mem_stage_inst_dmem_ram_154__10_), .C(mem_stage_inst_dmem_ram_153__10_), .D(mem_stage_inst_dmem_ram_155__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5194) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u564 ( .A(
        mem_stage_inst_dmem_ram_136__10_), .B(mem_stage_inst_dmem_ram_138__10_), .C(mem_stage_inst_dmem_ram_137__10_), .D(mem_stage_inst_dmem_ram_139__10_), 
        .S0(mem_stage_inst_dmem_n101), .S1(mem_stage_inst_dmem_n3), .Y(
        mem_stage_inst_dmem_n5199) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u563 ( .A(
        mem_stage_inst_dmem_ram_168__10_), .B(mem_stage_inst_dmem_ram_170__10_), .C(mem_stage_inst_dmem_ram_169__10_), .D(mem_stage_inst_dmem_ram_171__10_), 
        .S0(mem_stage_inst_dmem_n100), .S1(mem_stage_inst_dmem_n2), .Y(
        mem_stage_inst_dmem_n5189) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u562 ( .A(
        mem_stage_inst_dmem_ram_248__9_), .B(mem_stage_inst_dmem_ram_250__9_), 
        .C(mem_stage_inst_dmem_ram_249__9_), .D(
        mem_stage_inst_dmem_ram_251__9_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5080) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u561 ( .A(
        mem_stage_inst_dmem_ram_216__9_), .B(mem_stage_inst_dmem_ram_218__9_), 
        .C(mem_stage_inst_dmem_ram_217__9_), .D(
        mem_stage_inst_dmem_ram_219__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5090) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u560 ( .A(
        mem_stage_inst_dmem_ram_200__9_), .B(mem_stage_inst_dmem_ram_202__9_), 
        .C(mem_stage_inst_dmem_ram_201__9_), .D(
        mem_stage_inst_dmem_ram_203__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5095) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u559 ( .A(
        mem_stage_inst_dmem_ram_232__9_), .B(mem_stage_inst_dmem_ram_234__9_), 
        .C(mem_stage_inst_dmem_ram_233__9_), .D(
        mem_stage_inst_dmem_ram_235__9_), .S0(mem_stage_inst_dmem_n114), .S1(
        mem_stage_inst_dmem_n16), .Y(mem_stage_inst_dmem_n5085) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u558 ( .A(
        mem_stage_inst_dmem_ram_120__9_), .B(mem_stage_inst_dmem_ram_122__9_), 
        .C(mem_stage_inst_dmem_ram_121__9_), .D(
        mem_stage_inst_dmem_ram_123__9_), .S0(mem_stage_inst_dmem_n104), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5120) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u557 ( .A(mem_stage_inst_dmem_ram_88__9_), .B(mem_stage_inst_dmem_ram_90__9_), .C(mem_stage_inst_dmem_ram_89__9_), .D(
        mem_stage_inst_dmem_ram_91__9_), .S0(mem_stage_inst_dmem_n105), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5130) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u556 ( .A(mem_stage_inst_dmem_ram_72__9_), .B(mem_stage_inst_dmem_ram_74__9_), .C(mem_stage_inst_dmem_ram_73__9_), .D(
        mem_stage_inst_dmem_ram_75__9_), .S0(mem_stage_inst_dmem_n107), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n5135) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u555 ( .A(
        mem_stage_inst_dmem_ram_104__9_), .B(mem_stage_inst_dmem_ram_106__9_), 
        .C(mem_stage_inst_dmem_ram_105__9_), .D(
        mem_stage_inst_dmem_ram_107__9_), .S0(mem_stage_inst_dmem_n106), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5125) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u554 ( .A(mem_stage_inst_dmem_ram_56__9_), .B(mem_stage_inst_dmem_ram_58__9_), .C(mem_stage_inst_dmem_ram_57__9_), .D(
        mem_stage_inst_dmem_ram_59__9_), .S0(mem_stage_inst_dmem_n108), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n5140) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u553 ( .A(mem_stage_inst_dmem_ram_24__9_), .B(mem_stage_inst_dmem_ram_26__9_), .C(mem_stage_inst_dmem_ram_25__9_), .D(
        mem_stage_inst_dmem_ram_27__9_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n6), .Y(mem_stage_inst_dmem_n5150) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u552 ( .A(mem_stage_inst_dmem_ram_8__9_), 
        .B(mem_stage_inst_dmem_ram_10__9_), .C(mem_stage_inst_dmem_ram_9__9_), 
        .D(mem_stage_inst_dmem_ram_11__9_), .S0(mem_stage_inst_dmem_n121), 
        .S1(mem_stage_inst_dmem_n7), .Y(mem_stage_inst_dmem_n5155) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u551 ( .A(mem_stage_inst_dmem_ram_40__9_), .B(mem_stage_inst_dmem_ram_42__9_), .C(mem_stage_inst_dmem_ram_41__9_), .D(
        mem_stage_inst_dmem_ram_43__9_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n5145) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u550 ( .A(
        mem_stage_inst_dmem_ram_184__9_), .B(mem_stage_inst_dmem_ram_186__9_), 
        .C(mem_stage_inst_dmem_ram_185__9_), .D(
        mem_stage_inst_dmem_ram_187__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5100) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u549 ( .A(
        mem_stage_inst_dmem_ram_152__9_), .B(mem_stage_inst_dmem_ram_154__9_), 
        .C(mem_stage_inst_dmem_ram_153__9_), .D(
        mem_stage_inst_dmem_ram_155__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5110) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u548 ( .A(
        mem_stage_inst_dmem_ram_136__9_), .B(mem_stage_inst_dmem_ram_138__9_), 
        .C(mem_stage_inst_dmem_ram_137__9_), .D(
        mem_stage_inst_dmem_ram_139__9_), .S0(mem_stage_inst_dmem_n103), .S1(
        mem_stage_inst_dmem_n18), .Y(mem_stage_inst_dmem_n5115) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u547 ( .A(
        mem_stage_inst_dmem_ram_168__9_), .B(mem_stage_inst_dmem_ram_170__9_), 
        .C(mem_stage_inst_dmem_ram_169__9_), .D(
        mem_stage_inst_dmem_ram_171__9_), .S0(mem_stage_inst_dmem_n115), .S1(
        mem_stage_inst_dmem_n17), .Y(mem_stage_inst_dmem_n5105) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u546 ( .A(
        mem_stage_inst_dmem_ram_248__8_), .B(mem_stage_inst_dmem_ram_250__8_), 
        .C(mem_stage_inst_dmem_ram_249__8_), .D(
        mem_stage_inst_dmem_ram_251__8_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n4996) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u545 ( .A(
        mem_stage_inst_dmem_ram_216__8_), .B(mem_stage_inst_dmem_ram_218__8_), 
        .C(mem_stage_inst_dmem_ram_217__8_), .D(
        mem_stage_inst_dmem_ram_219__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5006) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u544 ( .A(
        mem_stage_inst_dmem_ram_200__8_), .B(mem_stage_inst_dmem_ram_202__8_), 
        .C(mem_stage_inst_dmem_ram_201__8_), .D(
        mem_stage_inst_dmem_ram_203__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5011) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u543 ( .A(
        mem_stage_inst_dmem_ram_232__8_), .B(mem_stage_inst_dmem_ram_234__8_), 
        .C(mem_stage_inst_dmem_ram_233__8_), .D(
        mem_stage_inst_dmem_ram_235__8_), .S0(mem_stage_inst_dmem_n109), .S1(
        mem_stage_inst_dmem_n11), .Y(mem_stage_inst_dmem_n5001) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u542 ( .A(
        mem_stage_inst_dmem_ram_120__8_), .B(mem_stage_inst_dmem_ram_122__8_), 
        .C(mem_stage_inst_dmem_ram_121__8_), .D(
        mem_stage_inst_dmem_ram_123__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5036) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u541 ( .A(mem_stage_inst_dmem_ram_88__8_), .B(mem_stage_inst_dmem_ram_90__8_), .C(mem_stage_inst_dmem_ram_89__8_), .D(
        mem_stage_inst_dmem_ram_91__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5046) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u540 ( .A(mem_stage_inst_dmem_ram_72__8_), .B(mem_stage_inst_dmem_ram_74__8_), .C(mem_stage_inst_dmem_ram_73__8_), .D(
        mem_stage_inst_dmem_ram_75__8_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5051) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u539 ( .A(
        mem_stage_inst_dmem_ram_104__8_), .B(mem_stage_inst_dmem_ram_106__8_), 
        .C(mem_stage_inst_dmem_ram_105__8_), .D(
        mem_stage_inst_dmem_ram_107__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5041) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u538 ( .A(mem_stage_inst_dmem_ram_56__8_), .B(mem_stage_inst_dmem_ram_58__8_), .C(mem_stage_inst_dmem_ram_57__8_), .D(
        mem_stage_inst_dmem_ram_59__8_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5056) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u537 ( .A(mem_stage_inst_dmem_ram_24__8_), .B(mem_stage_inst_dmem_ram_26__8_), .C(mem_stage_inst_dmem_ram_25__8_), .D(
        mem_stage_inst_dmem_ram_27__8_), .S0(mem_stage_inst_dmem_n113), .S1(
        mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5066) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u536 ( .A(mem_stage_inst_dmem_ram_8__8_), 
        .B(mem_stage_inst_dmem_ram_10__8_), .C(mem_stage_inst_dmem_ram_9__8_), 
        .D(mem_stage_inst_dmem_ram_11__8_), .S0(mem_stage_inst_dmem_n113), 
        .S1(mem_stage_inst_dmem_n15), .Y(mem_stage_inst_dmem_n5071) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u535 ( .A(mem_stage_inst_dmem_ram_40__8_), .B(mem_stage_inst_dmem_ram_42__8_), .C(mem_stage_inst_dmem_ram_41__8_), .D(
        mem_stage_inst_dmem_ram_43__8_), .S0(mem_stage_inst_dmem_n112), .S1(
        mem_stage_inst_dmem_n14), .Y(mem_stage_inst_dmem_n5061) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u534 ( .A(
        mem_stage_inst_dmem_ram_184__8_), .B(mem_stage_inst_dmem_ram_186__8_), 
        .C(mem_stage_inst_dmem_ram_185__8_), .D(
        mem_stage_inst_dmem_ram_187__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5016) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u533 ( .A(
        mem_stage_inst_dmem_ram_152__8_), .B(mem_stage_inst_dmem_ram_154__8_), 
        .C(mem_stage_inst_dmem_ram_153__8_), .D(
        mem_stage_inst_dmem_ram_155__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5026) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u532 ( .A(
        mem_stage_inst_dmem_ram_136__8_), .B(mem_stage_inst_dmem_ram_138__8_), 
        .C(mem_stage_inst_dmem_ram_137__8_), .D(
        mem_stage_inst_dmem_ram_139__8_), .S0(mem_stage_inst_dmem_n111), .S1(
        mem_stage_inst_dmem_n13), .Y(mem_stage_inst_dmem_n5031) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u531 ( .A(
        mem_stage_inst_dmem_ram_168__8_), .B(mem_stage_inst_dmem_ram_170__8_), 
        .C(mem_stage_inst_dmem_ram_169__8_), .D(
        mem_stage_inst_dmem_ram_171__8_), .S0(mem_stage_inst_dmem_n110), .S1(
        mem_stage_inst_dmem_n12), .Y(mem_stage_inst_dmem_n5021) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u530 ( .A(
        mem_stage_inst_dmem_ram_248__7_), .B(mem_stage_inst_dmem_ram_250__7_), 
        .C(mem_stage_inst_dmem_ram_249__7_), .D(
        mem_stage_inst_dmem_ram_251__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4912) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u529 ( .A(
        mem_stage_inst_dmem_ram_216__7_), .B(mem_stage_inst_dmem_ram_218__7_), 
        .C(mem_stage_inst_dmem_ram_217__7_), .D(
        mem_stage_inst_dmem_ram_219__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4922) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u528 ( .A(
        mem_stage_inst_dmem_ram_200__7_), .B(mem_stage_inst_dmem_ram_202__7_), 
        .C(mem_stage_inst_dmem_ram_201__7_), .D(
        mem_stage_inst_dmem_ram_203__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4927) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u527 ( .A(
        mem_stage_inst_dmem_ram_232__7_), .B(mem_stage_inst_dmem_ram_234__7_), 
        .C(mem_stage_inst_dmem_ram_233__7_), .D(
        mem_stage_inst_dmem_ram_235__7_), .S0(mem_stage_inst_dmem_n150), .S1(
        mem_stage_inst_dmem_n52), .Y(mem_stage_inst_dmem_n4917) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u526 ( .A(
        mem_stage_inst_dmem_ram_120__7_), .B(mem_stage_inst_dmem_ram_122__7_), 
        .C(mem_stage_inst_dmem_ram_121__7_), .D(
        mem_stage_inst_dmem_ram_123__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4952) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u525 ( .A(mem_stage_inst_dmem_ram_88__7_), .B(mem_stage_inst_dmem_ram_90__7_), .C(mem_stage_inst_dmem_ram_89__7_), .D(
        mem_stage_inst_dmem_ram_91__7_), .S0(mem_stage_inst_dmem_n153), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n4962) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u524 ( .A(mem_stage_inst_dmem_ram_72__7_), .B(mem_stage_inst_dmem_ram_74__7_), .C(mem_stage_inst_dmem_ram_73__7_), .D(
        mem_stage_inst_dmem_ram_75__7_), .S0(mem_stage_inst_dmem_n153), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n4967) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u523 ( .A(
        mem_stage_inst_dmem_ram_104__7_), .B(mem_stage_inst_dmem_ram_106__7_), 
        .C(mem_stage_inst_dmem_ram_105__7_), .D(
        mem_stage_inst_dmem_ram_107__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4957) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u522 ( .A(mem_stage_inst_dmem_ram_56__7_), .B(mem_stage_inst_dmem_ram_58__7_), .C(mem_stage_inst_dmem_ram_57__7_), .D(
        mem_stage_inst_dmem_ram_59__7_), .S0(mem_stage_inst_dmem_n153), .S1(
        mem_stage_inst_dmem_n55), .Y(mem_stage_inst_dmem_n4972) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u521 ( .A(mem_stage_inst_dmem_ram_24__7_), .B(mem_stage_inst_dmem_ram_26__7_), .C(mem_stage_inst_dmem_ram_25__7_), .D(
        mem_stage_inst_dmem_ram_27__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4982) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u520 ( .A(mem_stage_inst_dmem_ram_8__7_), 
        .B(mem_stage_inst_dmem_ram_10__7_), .C(mem_stage_inst_dmem_ram_9__7_), 
        .D(mem_stage_inst_dmem_ram_11__7_), .S0(mem_stage_inst_dmem_n154), 
        .S1(mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4987) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u519 ( .A(mem_stage_inst_dmem_ram_40__7_), .B(mem_stage_inst_dmem_ram_42__7_), .C(mem_stage_inst_dmem_ram_41__7_), .D(
        mem_stage_inst_dmem_ram_43__7_), .S0(mem_stage_inst_dmem_n154), .S1(
        mem_stage_inst_dmem_n56), .Y(mem_stage_inst_dmem_n4977) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u518 ( .A(
        mem_stage_inst_dmem_ram_184__7_), .B(mem_stage_inst_dmem_ram_186__7_), 
        .C(mem_stage_inst_dmem_ram_185__7_), .D(
        mem_stage_inst_dmem_ram_187__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4932) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u517 ( .A(
        mem_stage_inst_dmem_ram_152__7_), .B(mem_stage_inst_dmem_ram_154__7_), 
        .C(mem_stage_inst_dmem_ram_153__7_), .D(
        mem_stage_inst_dmem_ram_155__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4942) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u516 ( .A(
        mem_stage_inst_dmem_ram_136__7_), .B(mem_stage_inst_dmem_ram_138__7_), 
        .C(mem_stage_inst_dmem_ram_137__7_), .D(
        mem_stage_inst_dmem_ram_139__7_), .S0(mem_stage_inst_dmem_n152), .S1(
        mem_stage_inst_dmem_n54), .Y(mem_stage_inst_dmem_n4947) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u515 ( .A(
        mem_stage_inst_dmem_ram_168__7_), .B(mem_stage_inst_dmem_ram_170__7_), 
        .C(mem_stage_inst_dmem_ram_169__7_), .D(
        mem_stage_inst_dmem_ram_171__7_), .S0(mem_stage_inst_dmem_n151), .S1(
        mem_stage_inst_dmem_n53), .Y(mem_stage_inst_dmem_n4937) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u514 ( .A(
        mem_stage_inst_dmem_ram_248__6_), .B(mem_stage_inst_dmem_ram_250__6_), 
        .C(mem_stage_inst_dmem_ram_249__6_), .D(
        mem_stage_inst_dmem_ram_251__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4828) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u513 ( .A(
        mem_stage_inst_dmem_ram_216__6_), .B(mem_stage_inst_dmem_ram_218__6_), 
        .C(mem_stage_inst_dmem_ram_217__6_), .D(
        mem_stage_inst_dmem_ram_219__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4838) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u512 ( .A(
        mem_stage_inst_dmem_ram_200__6_), .B(mem_stage_inst_dmem_ram_202__6_), 
        .C(mem_stage_inst_dmem_ram_201__6_), .D(
        mem_stage_inst_dmem_ram_203__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4843) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u511 ( .A(
        mem_stage_inst_dmem_ram_232__6_), .B(mem_stage_inst_dmem_ram_234__6_), 
        .C(mem_stage_inst_dmem_ram_233__6_), .D(
        mem_stage_inst_dmem_ram_235__6_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n4833) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u510 ( .A(
        mem_stage_inst_dmem_ram_120__6_), .B(mem_stage_inst_dmem_ram_122__6_), 
        .C(mem_stage_inst_dmem_ram_121__6_), .D(
        mem_stage_inst_dmem_ram_123__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4868) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u509 ( .A(mem_stage_inst_dmem_ram_88__6_), .B(mem_stage_inst_dmem_ram_90__6_), .C(mem_stage_inst_dmem_ram_89__6_), .D(
        mem_stage_inst_dmem_ram_91__6_), .S0(mem_stage_inst_dmem_n148), .S1(
        mem_stage_inst_dmem_n50), .Y(mem_stage_inst_dmem_n4878) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u508 ( .A(mem_stage_inst_dmem_ram_72__6_), .B(mem_stage_inst_dmem_ram_74__6_), .C(mem_stage_inst_dmem_ram_73__6_), .D(
        mem_stage_inst_dmem_ram_75__6_), .S0(mem_stage_inst_dmem_n148), .S1(
        mem_stage_inst_dmem_n50), .Y(mem_stage_inst_dmem_n4883) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u507 ( .A(
        mem_stage_inst_dmem_ram_104__6_), .B(mem_stage_inst_dmem_ram_106__6_), 
        .C(mem_stage_inst_dmem_ram_105__6_), .D(
        mem_stage_inst_dmem_ram_107__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4873) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u506 ( .A(mem_stage_inst_dmem_ram_56__6_), .B(mem_stage_inst_dmem_ram_58__6_), .C(mem_stage_inst_dmem_ram_57__6_), .D(
        mem_stage_inst_dmem_ram_59__6_), .S0(mem_stage_inst_dmem_n148), .S1(
        mem_stage_inst_dmem_n50), .Y(mem_stage_inst_dmem_n4888) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u505 ( .A(mem_stage_inst_dmem_ram_24__6_), .B(mem_stage_inst_dmem_ram_26__6_), .C(mem_stage_inst_dmem_ram_25__6_), .D(
        mem_stage_inst_dmem_ram_27__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4898) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u504 ( .A(mem_stage_inst_dmem_ram_8__6_), 
        .B(mem_stage_inst_dmem_ram_10__6_), .C(mem_stage_inst_dmem_ram_9__6_), 
        .D(mem_stage_inst_dmem_ram_11__6_), .S0(mem_stage_inst_dmem_n149), 
        .S1(mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4903) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u503 ( .A(mem_stage_inst_dmem_ram_40__6_), .B(mem_stage_inst_dmem_ram_42__6_), .C(mem_stage_inst_dmem_ram_41__6_), .D(
        mem_stage_inst_dmem_ram_43__6_), .S0(mem_stage_inst_dmem_n149), .S1(
        mem_stage_inst_dmem_n51), .Y(mem_stage_inst_dmem_n4893) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u502 ( .A(
        mem_stage_inst_dmem_ram_184__6_), .B(mem_stage_inst_dmem_ram_186__6_), 
        .C(mem_stage_inst_dmem_ram_185__6_), .D(
        mem_stage_inst_dmem_ram_187__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4848) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u501 ( .A(
        mem_stage_inst_dmem_ram_152__6_), .B(mem_stage_inst_dmem_ram_154__6_), 
        .C(mem_stage_inst_dmem_ram_153__6_), .D(
        mem_stage_inst_dmem_ram_155__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4858) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u500 ( .A(
        mem_stage_inst_dmem_ram_136__6_), .B(mem_stage_inst_dmem_ram_138__6_), 
        .C(mem_stage_inst_dmem_ram_137__6_), .D(
        mem_stage_inst_dmem_ram_139__6_), .S0(mem_stage_inst_dmem_n147), .S1(
        mem_stage_inst_dmem_n49), .Y(mem_stage_inst_dmem_n4863) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u499 ( .A(
        mem_stage_inst_dmem_ram_168__6_), .B(mem_stage_inst_dmem_ram_170__6_), 
        .C(mem_stage_inst_dmem_ram_169__6_), .D(
        mem_stage_inst_dmem_ram_171__6_), .S0(mem_stage_inst_dmem_n146), .S1(
        mem_stage_inst_dmem_n48), .Y(mem_stage_inst_dmem_n4853) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u498 ( .A(
        mem_stage_inst_dmem_ram_248__5_), .B(mem_stage_inst_dmem_ram_250__5_), 
        .C(mem_stage_inst_dmem_ram_249__5_), .D(
        mem_stage_inst_dmem_ram_251__5_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4744) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u497 ( .A(
        mem_stage_inst_dmem_ram_216__5_), .B(mem_stage_inst_dmem_ram_218__5_), 
        .C(mem_stage_inst_dmem_ram_217__5_), .D(
        mem_stage_inst_dmem_ram_219__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4754) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u496 ( .A(
        mem_stage_inst_dmem_ram_200__5_), .B(mem_stage_inst_dmem_ram_202__5_), 
        .C(mem_stage_inst_dmem_ram_201__5_), .D(
        mem_stage_inst_dmem_ram_203__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4759) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u495 ( .A(
        mem_stage_inst_dmem_ram_232__5_), .B(mem_stage_inst_dmem_ram_234__5_), 
        .C(mem_stage_inst_dmem_ram_233__5_), .D(
        mem_stage_inst_dmem_ram_235__5_), .S0(mem_stage_inst_dmem_n160), .S1(
        mem_stage_inst_dmem_n62), .Y(mem_stage_inst_dmem_n4749) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u494 ( .A(
        mem_stage_inst_dmem_ram_120__5_), .B(mem_stage_inst_dmem_ram_122__5_), 
        .C(mem_stage_inst_dmem_ram_121__5_), .D(
        mem_stage_inst_dmem_ram_123__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4784) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u493 ( .A(mem_stage_inst_dmem_ram_88__5_), .B(mem_stage_inst_dmem_ram_90__5_), .C(mem_stage_inst_dmem_ram_89__5_), .D(
        mem_stage_inst_dmem_ram_91__5_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n4794) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u492 ( .A(mem_stage_inst_dmem_ram_72__5_), .B(mem_stage_inst_dmem_ram_74__5_), .C(mem_stage_inst_dmem_ram_73__5_), .D(
        mem_stage_inst_dmem_ram_75__5_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n4799) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u491 ( .A(
        mem_stage_inst_dmem_ram_104__5_), .B(mem_stage_inst_dmem_ram_106__5_), 
        .C(mem_stage_inst_dmem_ram_105__5_), .D(
        mem_stage_inst_dmem_ram_107__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4789) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u490 ( .A(mem_stage_inst_dmem_ram_56__5_), .B(mem_stage_inst_dmem_ram_58__5_), .C(mem_stage_inst_dmem_ram_57__5_), .D(
        mem_stage_inst_dmem_ram_59__5_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n4804) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u489 ( .A(mem_stage_inst_dmem_ram_24__5_), .B(mem_stage_inst_dmem_ram_26__5_), .C(mem_stage_inst_dmem_ram_25__5_), .D(
        mem_stage_inst_dmem_ram_27__5_), .S0(mem_stage_inst_dmem_n164), .S1(
        ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4814) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u488 ( .A(mem_stage_inst_dmem_ram_8__5_), 
        .B(mem_stage_inst_dmem_ram_10__5_), .C(mem_stage_inst_dmem_ram_9__5_), 
        .D(mem_stage_inst_dmem_ram_11__5_), .S0(mem_stage_inst_dmem_n164), 
        .S1(ex_pipeline_reg_out[22]), .Y(mem_stage_inst_dmem_n4819) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u487 ( .A(mem_stage_inst_dmem_ram_40__5_), .B(mem_stage_inst_dmem_ram_42__5_), .C(mem_stage_inst_dmem_ram_41__5_), .D(
        mem_stage_inst_dmem_ram_43__5_), .S0(mem_stage_inst_dmem_n163), .S1(
        mem_stage_inst_dmem_n65), .Y(mem_stage_inst_dmem_n4809) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u486 ( .A(
        mem_stage_inst_dmem_ram_184__5_), .B(mem_stage_inst_dmem_ram_186__5_), 
        .C(mem_stage_inst_dmem_ram_185__5_), .D(
        mem_stage_inst_dmem_ram_187__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4764) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u485 ( .A(
        mem_stage_inst_dmem_ram_152__5_), .B(mem_stage_inst_dmem_ram_154__5_), 
        .C(mem_stage_inst_dmem_ram_153__5_), .D(
        mem_stage_inst_dmem_ram_155__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4774) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u484 ( .A(
        mem_stage_inst_dmem_ram_136__5_), .B(mem_stage_inst_dmem_ram_138__5_), 
        .C(mem_stage_inst_dmem_ram_137__5_), .D(
        mem_stage_inst_dmem_ram_139__5_), .S0(mem_stage_inst_dmem_n162), .S1(
        mem_stage_inst_dmem_n64), .Y(mem_stage_inst_dmem_n4779) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u483 ( .A(
        mem_stage_inst_dmem_ram_168__5_), .B(mem_stage_inst_dmem_ram_170__5_), 
        .C(mem_stage_inst_dmem_ram_169__5_), .D(
        mem_stage_inst_dmem_ram_171__5_), .S0(mem_stage_inst_dmem_n161), .S1(
        mem_stage_inst_dmem_n63), .Y(mem_stage_inst_dmem_n4769) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u482 ( .A(
        mem_stage_inst_dmem_ram_248__4_), .B(mem_stage_inst_dmem_ram_250__4_), 
        .C(mem_stage_inst_dmem_ram_249__4_), .D(
        mem_stage_inst_dmem_ram_251__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n564) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u481 ( .A(
        mem_stage_inst_dmem_ram_216__4_), .B(mem_stage_inst_dmem_ram_218__4_), 
        .C(mem_stage_inst_dmem_ram_217__4_), .D(
        mem_stage_inst_dmem_ram_219__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4670) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u480 ( .A(
        mem_stage_inst_dmem_ram_200__4_), .B(mem_stage_inst_dmem_ram_202__4_), 
        .C(mem_stage_inst_dmem_ram_201__4_), .D(
        mem_stage_inst_dmem_ram_203__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4675) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u479 ( .A(
        mem_stage_inst_dmem_ram_232__4_), .B(mem_stage_inst_dmem_ram_234__4_), 
        .C(mem_stage_inst_dmem_ram_233__4_), .D(
        mem_stage_inst_dmem_ram_235__4_), .S0(mem_stage_inst_dmem_n155), .S1(
        mem_stage_inst_dmem_n57), .Y(mem_stage_inst_dmem_n4665) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u478 ( .A(
        mem_stage_inst_dmem_ram_120__4_), .B(mem_stage_inst_dmem_ram_122__4_), 
        .C(mem_stage_inst_dmem_ram_121__4_), .D(
        mem_stage_inst_dmem_ram_123__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4700) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u477 ( .A(mem_stage_inst_dmem_ram_88__4_), .B(mem_stage_inst_dmem_ram_90__4_), .C(mem_stage_inst_dmem_ram_89__4_), .D(
        mem_stage_inst_dmem_ram_91__4_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n4710) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u476 ( .A(mem_stage_inst_dmem_ram_72__4_), .B(mem_stage_inst_dmem_ram_74__4_), .C(mem_stage_inst_dmem_ram_73__4_), .D(
        mem_stage_inst_dmem_ram_75__4_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n4715) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u475 ( .A(
        mem_stage_inst_dmem_ram_104__4_), .B(mem_stage_inst_dmem_ram_106__4_), 
        .C(mem_stage_inst_dmem_ram_105__4_), .D(
        mem_stage_inst_dmem_ram_107__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4705) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u474 ( .A(mem_stage_inst_dmem_ram_56__4_), .B(mem_stage_inst_dmem_ram_58__4_), .C(mem_stage_inst_dmem_ram_57__4_), .D(
        mem_stage_inst_dmem_ram_59__4_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n4720) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u473 ( .A(mem_stage_inst_dmem_ram_24__4_), .B(mem_stage_inst_dmem_ram_26__4_), .C(mem_stage_inst_dmem_ram_25__4_), .D(
        mem_stage_inst_dmem_ram_27__4_), .S0(mem_stage_inst_dmem_n159), .S1(
        mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4730) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u472 ( .A(mem_stage_inst_dmem_ram_8__4_), 
        .B(mem_stage_inst_dmem_ram_10__4_), .C(mem_stage_inst_dmem_ram_9__4_), 
        .D(mem_stage_inst_dmem_ram_11__4_), .S0(mem_stage_inst_dmem_n159), 
        .S1(mem_stage_inst_dmem_n61), .Y(mem_stage_inst_dmem_n4735) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u471 ( .A(mem_stage_inst_dmem_ram_40__4_), .B(mem_stage_inst_dmem_ram_42__4_), .C(mem_stage_inst_dmem_ram_41__4_), .D(
        mem_stage_inst_dmem_ram_43__4_), .S0(mem_stage_inst_dmem_n158), .S1(
        mem_stage_inst_dmem_n60), .Y(mem_stage_inst_dmem_n4725) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u470 ( .A(
        mem_stage_inst_dmem_ram_184__4_), .B(mem_stage_inst_dmem_ram_186__4_), 
        .C(mem_stage_inst_dmem_ram_185__4_), .D(
        mem_stage_inst_dmem_ram_187__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4680) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u469 ( .A(
        mem_stage_inst_dmem_ram_152__4_), .B(mem_stage_inst_dmem_ram_154__4_), 
        .C(mem_stage_inst_dmem_ram_153__4_), .D(
        mem_stage_inst_dmem_ram_155__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4690) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u468 ( .A(
        mem_stage_inst_dmem_ram_136__4_), .B(mem_stage_inst_dmem_ram_138__4_), 
        .C(mem_stage_inst_dmem_ram_137__4_), .D(
        mem_stage_inst_dmem_ram_139__4_), .S0(mem_stage_inst_dmem_n157), .S1(
        mem_stage_inst_dmem_n59), .Y(mem_stage_inst_dmem_n4695) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u467 ( .A(
        mem_stage_inst_dmem_ram_168__4_), .B(mem_stage_inst_dmem_ram_170__4_), 
        .C(mem_stage_inst_dmem_ram_169__4_), .D(
        mem_stage_inst_dmem_ram_171__4_), .S0(mem_stage_inst_dmem_n156), .S1(
        mem_stage_inst_dmem_n58), .Y(mem_stage_inst_dmem_n4685) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u466 ( .A(
        mem_stage_inst_dmem_ram_248__3_), .B(mem_stage_inst_dmem_ram_250__3_), 
        .C(mem_stage_inst_dmem_ram_249__3_), .D(
        mem_stage_inst_dmem_ram_251__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n480) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u465 ( .A(
        mem_stage_inst_dmem_ram_216__3_), .B(mem_stage_inst_dmem_ram_218__3_), 
        .C(mem_stage_inst_dmem_ram_217__3_), .D(
        mem_stage_inst_dmem_ram_219__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n490) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u464 ( .A(
        mem_stage_inst_dmem_ram_200__3_), .B(mem_stage_inst_dmem_ram_202__3_), 
        .C(mem_stage_inst_dmem_ram_201__3_), .D(
        mem_stage_inst_dmem_ram_203__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n495) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u463 ( .A(
        mem_stage_inst_dmem_ram_232__3_), .B(mem_stage_inst_dmem_ram_234__3_), 
        .C(mem_stage_inst_dmem_ram_233__3_), .D(
        mem_stage_inst_dmem_ram_235__3_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n485) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u462 ( .A(
        mem_stage_inst_dmem_ram_120__3_), .B(mem_stage_inst_dmem_ram_122__3_), 
        .C(mem_stage_inst_dmem_ram_121__3_), .D(
        mem_stage_inst_dmem_ram_123__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n520) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u461 ( .A(mem_stage_inst_dmem_ram_88__3_), .B(mem_stage_inst_dmem_ram_90__3_), .C(mem_stage_inst_dmem_ram_89__3_), .D(
        mem_stage_inst_dmem_ram_91__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n530) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u460 ( .A(mem_stage_inst_dmem_ram_72__3_), .B(mem_stage_inst_dmem_ram_74__3_), .C(mem_stage_inst_dmem_ram_73__3_), .D(
        mem_stage_inst_dmem_ram_75__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n535) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u459 ( .A(
        mem_stage_inst_dmem_ram_104__3_), .B(mem_stage_inst_dmem_ram_106__3_), 
        .C(mem_stage_inst_dmem_ram_105__3_), .D(
        mem_stage_inst_dmem_ram_107__3_), .S0(mem_stage_inst_dmem_n133), .S1(
        mem_stage_inst_dmem_n35), .Y(mem_stage_inst_dmem_n525) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u458 ( .A(mem_stage_inst_dmem_ram_56__3_), .B(mem_stage_inst_dmem_ram_58__3_), .C(mem_stage_inst_dmem_ram_57__3_), .D(
        mem_stage_inst_dmem_ram_59__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n540) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u457 ( .A(mem_stage_inst_dmem_ram_24__3_), .B(mem_stage_inst_dmem_ram_26__3_), .C(mem_stage_inst_dmem_ram_25__3_), .D(
        mem_stage_inst_dmem_ram_27__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n550) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u456 ( .A(mem_stage_inst_dmem_ram_8__3_), 
        .B(mem_stage_inst_dmem_ram_10__3_), .C(mem_stage_inst_dmem_ram_9__3_), 
        .D(mem_stage_inst_dmem_ram_11__3_), .S0(mem_stage_inst_dmem_n135), 
        .S1(mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n555) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u455 ( .A(mem_stage_inst_dmem_ram_40__3_), .B(mem_stage_inst_dmem_ram_42__3_), .C(mem_stage_inst_dmem_ram_41__3_), .D(
        mem_stage_inst_dmem_ram_43__3_), .S0(mem_stage_inst_dmem_n134), .S1(
        mem_stage_inst_dmem_n36), .Y(mem_stage_inst_dmem_n545) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u454 ( .A(
        mem_stage_inst_dmem_ram_184__3_), .B(mem_stage_inst_dmem_ram_186__3_), 
        .C(mem_stage_inst_dmem_ram_185__3_), .D(
        mem_stage_inst_dmem_ram_187__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n500) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u453 ( .A(
        mem_stage_inst_dmem_ram_152__3_), .B(mem_stage_inst_dmem_ram_154__3_), 
        .C(mem_stage_inst_dmem_ram_153__3_), .D(
        mem_stage_inst_dmem_ram_155__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n510) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u452 ( .A(
        mem_stage_inst_dmem_ram_136__3_), .B(mem_stage_inst_dmem_ram_138__3_), 
        .C(mem_stage_inst_dmem_ram_137__3_), .D(
        mem_stage_inst_dmem_ram_139__3_), .S0(mem_stage_inst_dmem_n132), .S1(
        mem_stage_inst_dmem_n34), .Y(mem_stage_inst_dmem_n515) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u451 ( .A(
        mem_stage_inst_dmem_ram_168__3_), .B(mem_stage_inst_dmem_ram_170__3_), 
        .C(mem_stage_inst_dmem_ram_169__3_), .D(
        mem_stage_inst_dmem_ram_171__3_), .S0(mem_stage_inst_dmem_n131), .S1(
        mem_stage_inst_dmem_n33), .Y(mem_stage_inst_dmem_n505) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u450 ( .A(
        mem_stage_inst_dmem_ram_248__2_), .B(mem_stage_inst_dmem_ram_250__2_), 
        .C(mem_stage_inst_dmem_ram_249__2_), .D(
        mem_stage_inst_dmem_ram_251__2_), .S0(mem_stage_inst_dmem_n130), .S1(
        mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n396) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u449 ( .A(
        mem_stage_inst_dmem_ram_216__2_), .B(mem_stage_inst_dmem_ram_218__2_), 
        .C(mem_stage_inst_dmem_ram_217__2_), .D(
        mem_stage_inst_dmem_ram_219__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n406) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u448 ( .A(
        mem_stage_inst_dmem_ram_200__2_), .B(mem_stage_inst_dmem_ram_202__2_), 
        .C(mem_stage_inst_dmem_ram_201__2_), .D(
        mem_stage_inst_dmem_ram_203__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n411) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u447 ( .A(
        mem_stage_inst_dmem_ram_232__2_), .B(mem_stage_inst_dmem_ram_234__2_), 
        .C(mem_stage_inst_dmem_ram_233__2_), .D(
        mem_stage_inst_dmem_ram_235__2_), .S0(mem_stage_inst_dmem_n125), .S1(
        mem_stage_inst_dmem_n27), .Y(mem_stage_inst_dmem_n401) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u446 ( .A(
        mem_stage_inst_dmem_ram_120__2_), .B(mem_stage_inst_dmem_ram_122__2_), 
        .C(mem_stage_inst_dmem_ram_121__2_), .D(
        mem_stage_inst_dmem_ram_123__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n436) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u445 ( .A(mem_stage_inst_dmem_ram_88__2_), .B(mem_stage_inst_dmem_ram_90__2_), .C(mem_stage_inst_dmem_ram_89__2_), .D(
        mem_stage_inst_dmem_ram_91__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n446) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u444 ( .A(mem_stage_inst_dmem_ram_72__2_), .B(mem_stage_inst_dmem_ram_74__2_), .C(mem_stage_inst_dmem_ram_73__2_), .D(
        mem_stage_inst_dmem_ram_75__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n451) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u443 ( .A(
        mem_stage_inst_dmem_ram_104__2_), .B(mem_stage_inst_dmem_ram_106__2_), 
        .C(mem_stage_inst_dmem_ram_105__2_), .D(
        mem_stage_inst_dmem_ram_107__2_), .S0(mem_stage_inst_dmem_n128), .S1(
        mem_stage_inst_dmem_n30), .Y(mem_stage_inst_dmem_n441) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u442 ( .A(mem_stage_inst_dmem_ram_56__2_), .B(mem_stage_inst_dmem_ram_58__2_), .C(mem_stage_inst_dmem_ram_57__2_), .D(
        mem_stage_inst_dmem_ram_59__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n456) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u441 ( .A(mem_stage_inst_dmem_ram_24__2_), .B(mem_stage_inst_dmem_ram_26__2_), .C(mem_stage_inst_dmem_ram_25__2_), .D(
        mem_stage_inst_dmem_ram_27__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n466) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u440 ( .A(mem_stage_inst_dmem_ram_8__2_), 
        .B(mem_stage_inst_dmem_ram_10__2_), .C(mem_stage_inst_dmem_ram_9__2_), 
        .D(mem_stage_inst_dmem_ram_11__2_), .S0(mem_stage_inst_dmem_n130), 
        .S1(mem_stage_inst_dmem_n32), .Y(mem_stage_inst_dmem_n471) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u439 ( .A(mem_stage_inst_dmem_ram_40__2_), .B(mem_stage_inst_dmem_ram_42__2_), .C(mem_stage_inst_dmem_ram_41__2_), .D(
        mem_stage_inst_dmem_ram_43__2_), .S0(mem_stage_inst_dmem_n129), .S1(
        mem_stage_inst_dmem_n31), .Y(mem_stage_inst_dmem_n461) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u438 ( .A(
        mem_stage_inst_dmem_ram_184__2_), .B(mem_stage_inst_dmem_ram_186__2_), 
        .C(mem_stage_inst_dmem_ram_185__2_), .D(
        mem_stage_inst_dmem_ram_187__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n416) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u437 ( .A(
        mem_stage_inst_dmem_ram_152__2_), .B(mem_stage_inst_dmem_ram_154__2_), 
        .C(mem_stage_inst_dmem_ram_153__2_), .D(
        mem_stage_inst_dmem_ram_155__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n426) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u436 ( .A(
        mem_stage_inst_dmem_ram_136__2_), .B(mem_stage_inst_dmem_ram_138__2_), 
        .C(mem_stage_inst_dmem_ram_137__2_), .D(
        mem_stage_inst_dmem_ram_139__2_), .S0(mem_stage_inst_dmem_n127), .S1(
        mem_stage_inst_dmem_n29), .Y(mem_stage_inst_dmem_n431) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u435 ( .A(
        mem_stage_inst_dmem_ram_168__2_), .B(mem_stage_inst_dmem_ram_170__2_), 
        .C(mem_stage_inst_dmem_ram_169__2_), .D(
        mem_stage_inst_dmem_ram_171__2_), .S0(mem_stage_inst_dmem_n126), .S1(
        mem_stage_inst_dmem_n28), .Y(mem_stage_inst_dmem_n421) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u434 ( .A(
        mem_stage_inst_dmem_ram_248__1_), .B(mem_stage_inst_dmem_ram_250__1_), 
        .C(mem_stage_inst_dmem_ram_249__1_), .D(
        mem_stage_inst_dmem_ram_251__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n312) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u433 ( .A(
        mem_stage_inst_dmem_ram_216__1_), .B(mem_stage_inst_dmem_ram_218__1_), 
        .C(mem_stage_inst_dmem_ram_217__1_), .D(
        mem_stage_inst_dmem_ram_219__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n322) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u432 ( .A(
        mem_stage_inst_dmem_ram_200__1_), .B(mem_stage_inst_dmem_ram_202__1_), 
        .C(mem_stage_inst_dmem_ram_201__1_), .D(
        mem_stage_inst_dmem_ram_203__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n327) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u431 ( .A(
        mem_stage_inst_dmem_ram_232__1_), .B(mem_stage_inst_dmem_ram_234__1_), 
        .C(mem_stage_inst_dmem_ram_233__1_), .D(
        mem_stage_inst_dmem_ram_235__1_), .S0(mem_stage_inst_dmem_n140), .S1(
        mem_stage_inst_dmem_n42), .Y(mem_stage_inst_dmem_n317) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u430 ( .A(
        mem_stage_inst_dmem_ram_120__1_), .B(mem_stage_inst_dmem_ram_122__1_), 
        .C(mem_stage_inst_dmem_ram_121__1_), .D(
        mem_stage_inst_dmem_ram_123__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n352) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u429 ( .A(mem_stage_inst_dmem_ram_88__1_), .B(mem_stage_inst_dmem_ram_90__1_), .C(mem_stage_inst_dmem_ram_89__1_), .D(
        mem_stage_inst_dmem_ram_91__1_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n362) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u428 ( .A(mem_stage_inst_dmem_ram_72__1_), .B(mem_stage_inst_dmem_ram_74__1_), .C(mem_stage_inst_dmem_ram_73__1_), .D(
        mem_stage_inst_dmem_ram_75__1_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n367) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u427 ( .A(
        mem_stage_inst_dmem_ram_104__1_), .B(mem_stage_inst_dmem_ram_106__1_), 
        .C(mem_stage_inst_dmem_ram_105__1_), .D(
        mem_stage_inst_dmem_ram_107__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n357) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u426 ( .A(mem_stage_inst_dmem_ram_56__1_), .B(mem_stage_inst_dmem_ram_58__1_), .C(mem_stage_inst_dmem_ram_57__1_), .D(
        mem_stage_inst_dmem_ram_59__1_), .S0(mem_stage_inst_dmem_n143), .S1(
        mem_stage_inst_dmem_n45), .Y(mem_stage_inst_dmem_n372) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u425 ( .A(mem_stage_inst_dmem_ram_24__1_), .B(mem_stage_inst_dmem_ram_26__1_), .C(mem_stage_inst_dmem_ram_25__1_), .D(
        mem_stage_inst_dmem_ram_27__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n382) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u424 ( .A(mem_stage_inst_dmem_ram_8__1_), 
        .B(mem_stage_inst_dmem_ram_10__1_), .C(mem_stage_inst_dmem_ram_9__1_), 
        .D(mem_stage_inst_dmem_ram_11__1_), .S0(mem_stage_inst_dmem_n144), 
        .S1(mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n387) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u423 ( .A(mem_stage_inst_dmem_ram_40__1_), .B(mem_stage_inst_dmem_ram_42__1_), .C(mem_stage_inst_dmem_ram_41__1_), .D(
        mem_stage_inst_dmem_ram_43__1_), .S0(mem_stage_inst_dmem_n144), .S1(
        mem_stage_inst_dmem_n46), .Y(mem_stage_inst_dmem_n377) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u422 ( .A(
        mem_stage_inst_dmem_ram_184__1_), .B(mem_stage_inst_dmem_ram_186__1_), 
        .C(mem_stage_inst_dmem_ram_185__1_), .D(
        mem_stage_inst_dmem_ram_187__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n332) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u421 ( .A(
        mem_stage_inst_dmem_ram_152__1_), .B(mem_stage_inst_dmem_ram_154__1_), 
        .C(mem_stage_inst_dmem_ram_153__1_), .D(
        mem_stage_inst_dmem_ram_155__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n342) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u420 ( .A(
        mem_stage_inst_dmem_ram_136__1_), .B(mem_stage_inst_dmem_ram_138__1_), 
        .C(mem_stage_inst_dmem_ram_137__1_), .D(
        mem_stage_inst_dmem_ram_139__1_), .S0(mem_stage_inst_dmem_n142), .S1(
        mem_stage_inst_dmem_n44), .Y(mem_stage_inst_dmem_n347) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u419 ( .A(
        mem_stage_inst_dmem_ram_168__1_), .B(mem_stage_inst_dmem_ram_170__1_), 
        .C(mem_stage_inst_dmem_ram_169__1_), .D(
        mem_stage_inst_dmem_ram_171__1_), .S0(mem_stage_inst_dmem_n141), .S1(
        mem_stage_inst_dmem_n43), .Y(mem_stage_inst_dmem_n337) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u418 ( .A(
        mem_stage_inst_dmem_ram_248__0_), .B(mem_stage_inst_dmem_ram_250__0_), 
        .C(mem_stage_inst_dmem_ram_249__0_), .D(
        mem_stage_inst_dmem_ram_251__0_), .S0(mem_stage_inst_dmem_n145), .S1(
        mem_stage_inst_dmem_n47), .Y(mem_stage_inst_dmem_n228) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u417 ( .A(
        mem_stage_inst_dmem_ram_216__0_), .B(mem_stage_inst_dmem_ram_218__0_), 
        .C(mem_stage_inst_dmem_ram_217__0_), .D(
        mem_stage_inst_dmem_ram_219__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n238) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u416 ( .A(
        mem_stage_inst_dmem_ram_200__0_), .B(mem_stage_inst_dmem_ram_202__0_), 
        .C(mem_stage_inst_dmem_ram_201__0_), .D(
        mem_stage_inst_dmem_ram_203__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n243) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u415 ( .A(
        mem_stage_inst_dmem_ram_232__0_), .B(mem_stage_inst_dmem_ram_234__0_), 
        .C(mem_stage_inst_dmem_ram_233__0_), .D(
        mem_stage_inst_dmem_ram_235__0_), .S0(mem_stage_inst_dmem_n135), .S1(
        mem_stage_inst_dmem_n37), .Y(mem_stage_inst_dmem_n233) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u414 ( .A(
        mem_stage_inst_dmem_ram_120__0_), .B(mem_stage_inst_dmem_ram_122__0_), 
        .C(mem_stage_inst_dmem_ram_121__0_), .D(
        mem_stage_inst_dmem_ram_123__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n268) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u413 ( .A(mem_stage_inst_dmem_ram_88__0_), .B(mem_stage_inst_dmem_ram_90__0_), .C(mem_stage_inst_dmem_ram_89__0_), .D(
        mem_stage_inst_dmem_ram_91__0_), .S0(mem_stage_inst_dmem_n138), .S1(
        mem_stage_inst_dmem_n40), .Y(mem_stage_inst_dmem_n278) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u412 ( .A(mem_stage_inst_dmem_ram_72__0_), .B(mem_stage_inst_dmem_ram_74__0_), .C(mem_stage_inst_dmem_ram_73__0_), .D(
        mem_stage_inst_dmem_ram_75__0_), .S0(mem_stage_inst_dmem_n138), .S1(
        mem_stage_inst_dmem_n40), .Y(mem_stage_inst_dmem_n283) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u411 ( .A(
        mem_stage_inst_dmem_ram_104__0_), .B(mem_stage_inst_dmem_ram_106__0_), 
        .C(mem_stage_inst_dmem_ram_105__0_), .D(
        mem_stage_inst_dmem_ram_107__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n273) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u410 ( .A(mem_stage_inst_dmem_ram_56__0_), .B(mem_stage_inst_dmem_ram_58__0_), .C(mem_stage_inst_dmem_ram_57__0_), .D(
        mem_stage_inst_dmem_ram_59__0_), .S0(mem_stage_inst_dmem_n138), .S1(
        mem_stage_inst_dmem_n40), .Y(mem_stage_inst_dmem_n288) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u409 ( .A(mem_stage_inst_dmem_ram_24__0_), .B(mem_stage_inst_dmem_ram_26__0_), .C(mem_stage_inst_dmem_ram_25__0_), .D(
        mem_stage_inst_dmem_ram_27__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n298) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u408 ( .A(mem_stage_inst_dmem_ram_8__0_), 
        .B(mem_stage_inst_dmem_ram_10__0_), .C(mem_stage_inst_dmem_ram_9__0_), 
        .D(mem_stage_inst_dmem_ram_11__0_), .S0(mem_stage_inst_dmem_n139), 
        .S1(mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n303) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u407 ( .A(mem_stage_inst_dmem_ram_40__0_), .B(mem_stage_inst_dmem_ram_42__0_), .C(mem_stage_inst_dmem_ram_41__0_), .D(
        mem_stage_inst_dmem_ram_43__0_), .S0(mem_stage_inst_dmem_n139), .S1(
        mem_stage_inst_dmem_n41), .Y(mem_stage_inst_dmem_n293) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u406 ( .A(
        mem_stage_inst_dmem_ram_184__0_), .B(mem_stage_inst_dmem_ram_186__0_), 
        .C(mem_stage_inst_dmem_ram_185__0_), .D(
        mem_stage_inst_dmem_ram_187__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n248) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u405 ( .A(
        mem_stage_inst_dmem_ram_152__0_), .B(mem_stage_inst_dmem_ram_154__0_), 
        .C(mem_stage_inst_dmem_ram_153__0_), .D(
        mem_stage_inst_dmem_ram_155__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n258) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u404 ( .A(
        mem_stage_inst_dmem_ram_136__0_), .B(mem_stage_inst_dmem_ram_138__0_), 
        .C(mem_stage_inst_dmem_ram_137__0_), .D(
        mem_stage_inst_dmem_ram_139__0_), .S0(mem_stage_inst_dmem_n137), .S1(
        mem_stage_inst_dmem_n39), .Y(mem_stage_inst_dmem_n263) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u403 ( .A(
        mem_stage_inst_dmem_ram_168__0_), .B(mem_stage_inst_dmem_ram_170__0_), 
        .C(mem_stage_inst_dmem_ram_169__0_), .D(
        mem_stage_inst_dmem_ram_171__0_), .S0(mem_stage_inst_dmem_n136), .S1(
        mem_stage_inst_dmem_n38), .Y(mem_stage_inst_dmem_n253) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u402 ( .A(mem_stage_inst_dmem_n5658), 
        .B(mem_stage_inst_dmem_n5659), .C(mem_stage_inst_dmem_n5660), .D(
        mem_stage_inst_dmem_n5661), .S0(mem_stage_inst_dmem_n212), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5657) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u401 ( .A(mem_stage_inst_dmem_n5653), 
        .B(mem_stage_inst_dmem_n5654), .C(mem_stage_inst_dmem_n5655), .D(
        mem_stage_inst_dmem_n5656), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5652) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u400 ( .A(mem_stage_inst_dmem_n5643), 
        .B(mem_stage_inst_dmem_n5644), .C(mem_stage_inst_dmem_n5645), .D(
        mem_stage_inst_dmem_n5646), .S0(ex_pipeline_reg_out[25]), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5642) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u399 ( .A(mem_stage_inst_dmem_n5657), 
        .B(mem_stage_inst_dmem_n5647), .C(mem_stage_inst_dmem_n5652), .D(
        mem_stage_inst_dmem_n5642), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5662) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u398 ( .A(mem_stage_inst_dmem_n5574), 
        .B(mem_stage_inst_dmem_n5575), .C(mem_stage_inst_dmem_n5576), .D(
        mem_stage_inst_dmem_n5577), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5573) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u397 ( .A(mem_stage_inst_dmem_n5569), 
        .B(mem_stage_inst_dmem_n5570), .C(mem_stage_inst_dmem_n5571), .D(
        mem_stage_inst_dmem_n5572), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5568) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u396 ( .A(mem_stage_inst_dmem_n5559), 
        .B(mem_stage_inst_dmem_n5560), .C(mem_stage_inst_dmem_n5561), .D(
        mem_stage_inst_dmem_n5562), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5558) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u395 ( .A(mem_stage_inst_dmem_n5573), 
        .B(mem_stage_inst_dmem_n5563), .C(mem_stage_inst_dmem_n5568), .D(
        mem_stage_inst_dmem_n5558), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5578) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u394 ( .A(mem_stage_inst_dmem_n5490), 
        .B(mem_stage_inst_dmem_n5491), .C(mem_stage_inst_dmem_n5492), .D(
        mem_stage_inst_dmem_n5493), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5489) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u393 ( .A(mem_stage_inst_dmem_n5485), 
        .B(mem_stage_inst_dmem_n5486), .C(mem_stage_inst_dmem_n5487), .D(
        mem_stage_inst_dmem_n5488), .S0(mem_stage_inst_dmem_n212), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5484) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u392 ( .A(mem_stage_inst_dmem_n5475), 
        .B(mem_stage_inst_dmem_n5476), .C(mem_stage_inst_dmem_n5477), .D(
        mem_stage_inst_dmem_n5478), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5474) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u391 ( .A(mem_stage_inst_dmem_n5489), 
        .B(mem_stage_inst_dmem_n5479), .C(mem_stage_inst_dmem_n5484), .D(
        mem_stage_inst_dmem_n5474), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5494) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u390 ( .A(mem_stage_inst_dmem_n5406), 
        .B(mem_stage_inst_dmem_n5407), .C(mem_stage_inst_dmem_n5408), .D(
        mem_stage_inst_dmem_n5409), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5405) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u389 ( .A(mem_stage_inst_dmem_n5401), 
        .B(mem_stage_inst_dmem_n5402), .C(mem_stage_inst_dmem_n5403), .D(
        mem_stage_inst_dmem_n5404), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5400) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u388 ( .A(mem_stage_inst_dmem_n5391), 
        .B(mem_stage_inst_dmem_n5392), .C(mem_stage_inst_dmem_n5393), .D(
        mem_stage_inst_dmem_n5394), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5390) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u387 ( .A(mem_stage_inst_dmem_n5405), 
        .B(mem_stage_inst_dmem_n5395), .C(mem_stage_inst_dmem_n5400), .D(
        mem_stage_inst_dmem_n5390), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5410) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u386 ( .A(mem_stage_inst_dmem_n5322), 
        .B(mem_stage_inst_dmem_n5323), .C(mem_stage_inst_dmem_n5324), .D(
        mem_stage_inst_dmem_n5325), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5321) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u385 ( .A(mem_stage_inst_dmem_n5317), 
        .B(mem_stage_inst_dmem_n5318), .C(mem_stage_inst_dmem_n5319), .D(
        mem_stage_inst_dmem_n5320), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5316) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u384 ( .A(mem_stage_inst_dmem_n5307), 
        .B(mem_stage_inst_dmem_n5308), .C(mem_stage_inst_dmem_n5309), .D(
        mem_stage_inst_dmem_n5310), .S0(mem_stage_inst_dmem_n216), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5306) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u383 ( .A(mem_stage_inst_dmem_n5321), 
        .B(mem_stage_inst_dmem_n5311), .C(mem_stage_inst_dmem_n5316), .D(
        mem_stage_inst_dmem_n5306), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5326) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u382 ( .A(mem_stage_inst_dmem_n5238), 
        .B(mem_stage_inst_dmem_n5239), .C(mem_stage_inst_dmem_n5240), .D(
        mem_stage_inst_dmem_n5241), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5237) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u381 ( .A(mem_stage_inst_dmem_n5233), 
        .B(mem_stage_inst_dmem_n5234), .C(mem_stage_inst_dmem_n5235), .D(
        mem_stage_inst_dmem_n5236), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5232) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u380 ( .A(mem_stage_inst_dmem_n5223), 
        .B(mem_stage_inst_dmem_n5224), .C(mem_stage_inst_dmem_n5225), .D(
        mem_stage_inst_dmem_n5226), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5222) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u379 ( .A(mem_stage_inst_dmem_n5237), 
        .B(mem_stage_inst_dmem_n5227), .C(mem_stage_inst_dmem_n5232), .D(
        mem_stage_inst_dmem_n5222), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5242) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u378 ( .A(mem_stage_inst_dmem_n5154), 
        .B(mem_stage_inst_dmem_n5155), .C(mem_stage_inst_dmem_n5156), .D(
        mem_stage_inst_dmem_n5157), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5153) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u377 ( .A(mem_stage_inst_dmem_n5149), 
        .B(mem_stage_inst_dmem_n5150), .C(mem_stage_inst_dmem_n5151), .D(
        mem_stage_inst_dmem_n5152), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5148) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u376 ( .A(mem_stage_inst_dmem_n5139), 
        .B(mem_stage_inst_dmem_n5140), .C(mem_stage_inst_dmem_n5141), .D(
        mem_stage_inst_dmem_n5142), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5138) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u375 ( .A(mem_stage_inst_dmem_n5153), 
        .B(mem_stage_inst_dmem_n5143), .C(mem_stage_inst_dmem_n5148), .D(
        mem_stage_inst_dmem_n5138), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5158) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u374 ( .A(mem_stage_inst_dmem_n5070), 
        .B(mem_stage_inst_dmem_n5071), .C(mem_stage_inst_dmem_n5072), .D(
        mem_stage_inst_dmem_n5073), .S0(mem_stage_inst_dmem_n214), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5069) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u373 ( .A(mem_stage_inst_dmem_n5065), 
        .B(mem_stage_inst_dmem_n5066), .C(mem_stage_inst_dmem_n5067), .D(
        mem_stage_inst_dmem_n5068), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5064) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u372 ( .A(mem_stage_inst_dmem_n5055), 
        .B(mem_stage_inst_dmem_n5056), .C(mem_stage_inst_dmem_n5057), .D(
        mem_stage_inst_dmem_n5058), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5054) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u371 ( .A(mem_stage_inst_dmem_n5069), 
        .B(mem_stage_inst_dmem_n5059), .C(mem_stage_inst_dmem_n5064), .D(
        mem_stage_inst_dmem_n5054), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5074) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u370 ( .A(mem_stage_inst_dmem_n4986), 
        .B(mem_stage_inst_dmem_n4987), .C(mem_stage_inst_dmem_n4988), .D(
        mem_stage_inst_dmem_n4989), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4985) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u369 ( .A(mem_stage_inst_dmem_n4981), 
        .B(mem_stage_inst_dmem_n4982), .C(mem_stage_inst_dmem_n4983), .D(
        mem_stage_inst_dmem_n4984), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4980) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u368 ( .A(mem_stage_inst_dmem_n4971), 
        .B(mem_stage_inst_dmem_n4972), .C(mem_stage_inst_dmem_n4973), .D(
        mem_stage_inst_dmem_n4974), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4970) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u367 ( .A(mem_stage_inst_dmem_n4985), 
        .B(mem_stage_inst_dmem_n4975), .C(mem_stage_inst_dmem_n4980), .D(
        mem_stage_inst_dmem_n4970), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4990) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u366 ( .A(mem_stage_inst_dmem_n4902), 
        .B(mem_stage_inst_dmem_n4903), .C(mem_stage_inst_dmem_n4904), .D(
        mem_stage_inst_dmem_n4905), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4901) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u365 ( .A(mem_stage_inst_dmem_n4897), 
        .B(mem_stage_inst_dmem_n4898), .C(mem_stage_inst_dmem_n4899), .D(
        mem_stage_inst_dmem_n4900), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4896) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u364 ( .A(mem_stage_inst_dmem_n4887), 
        .B(mem_stage_inst_dmem_n4888), .C(mem_stage_inst_dmem_n4889), .D(
        mem_stage_inst_dmem_n4890), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4886) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u363 ( .A(mem_stage_inst_dmem_n4901), 
        .B(mem_stage_inst_dmem_n4891), .C(mem_stage_inst_dmem_n4896), .D(
        mem_stage_inst_dmem_n4886), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4906) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u362 ( .A(mem_stage_inst_dmem_n4818), 
        .B(mem_stage_inst_dmem_n4819), .C(mem_stage_inst_dmem_n4820), .D(
        mem_stage_inst_dmem_n4821), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4817) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u361 ( .A(mem_stage_inst_dmem_n4813), 
        .B(mem_stage_inst_dmem_n4814), .C(mem_stage_inst_dmem_n4815), .D(
        mem_stage_inst_dmem_n4816), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4812) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u360 ( .A(mem_stage_inst_dmem_n4803), 
        .B(mem_stage_inst_dmem_n4804), .C(mem_stage_inst_dmem_n4805), .D(
        mem_stage_inst_dmem_n4806), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4802) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u359 ( .A(mem_stage_inst_dmem_n4817), 
        .B(mem_stage_inst_dmem_n4807), .C(mem_stage_inst_dmem_n4812), .D(
        mem_stage_inst_dmem_n4802), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4822) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u358 ( .A(mem_stage_inst_dmem_n4734), 
        .B(mem_stage_inst_dmem_n4735), .C(mem_stage_inst_dmem_n4736), .D(
        mem_stage_inst_dmem_n4737), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4733) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u357 ( .A(mem_stage_inst_dmem_n4729), 
        .B(mem_stage_inst_dmem_n4730), .C(mem_stage_inst_dmem_n4731), .D(
        mem_stage_inst_dmem_n4732), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4728) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u356 ( .A(mem_stage_inst_dmem_n4719), 
        .B(mem_stage_inst_dmem_n4720), .C(mem_stage_inst_dmem_n4721), .D(
        mem_stage_inst_dmem_n4722), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4718) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u355 ( .A(mem_stage_inst_dmem_n4733), 
        .B(mem_stage_inst_dmem_n4723), .C(mem_stage_inst_dmem_n4728), .D(
        mem_stage_inst_dmem_n4718), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4738) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u354 ( .A(mem_stage_inst_dmem_n554), .B(
        mem_stage_inst_dmem_n555), .C(mem_stage_inst_dmem_n556), .D(
        mem_stage_inst_dmem_n557), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n553) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u353 ( .A(mem_stage_inst_dmem_n549), .B(
        mem_stage_inst_dmem_n550), .C(mem_stage_inst_dmem_n551), .D(
        mem_stage_inst_dmem_n552), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n548) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u352 ( .A(mem_stage_inst_dmem_n539), .B(
        mem_stage_inst_dmem_n540), .C(mem_stage_inst_dmem_n541), .D(
        mem_stage_inst_dmem_n542), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n538) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u351 ( .A(mem_stage_inst_dmem_n553), .B(
        mem_stage_inst_dmem_n543), .C(mem_stage_inst_dmem_n548), .D(
        mem_stage_inst_dmem_n538), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n558) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u350 ( .A(mem_stage_inst_dmem_n470), .B(
        mem_stage_inst_dmem_n471), .C(mem_stage_inst_dmem_n472), .D(
        mem_stage_inst_dmem_n473), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n469) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u349 ( .A(mem_stage_inst_dmem_n465), .B(
        mem_stage_inst_dmem_n466), .C(mem_stage_inst_dmem_n467), .D(
        mem_stage_inst_dmem_n468), .S0(mem_stage_inst_dmem_n210), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n464) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u348 ( .A(mem_stage_inst_dmem_n455), .B(
        mem_stage_inst_dmem_n456), .C(mem_stage_inst_dmem_n457), .D(
        mem_stage_inst_dmem_n458), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n454) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u347 ( .A(mem_stage_inst_dmem_n469), .B(
        mem_stage_inst_dmem_n459), .C(mem_stage_inst_dmem_n464), .D(
        mem_stage_inst_dmem_n454), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n474) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u346 ( .A(mem_stage_inst_dmem_n386), .B(
        mem_stage_inst_dmem_n387), .C(mem_stage_inst_dmem_n388), .D(
        mem_stage_inst_dmem_n389), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n385) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u345 ( .A(mem_stage_inst_dmem_n381), .B(
        mem_stage_inst_dmem_n382), .C(mem_stage_inst_dmem_n383), .D(
        mem_stage_inst_dmem_n384), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n380) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u344 ( .A(mem_stage_inst_dmem_n371), .B(
        mem_stage_inst_dmem_n372), .C(mem_stage_inst_dmem_n373), .D(
        mem_stage_inst_dmem_n374), .S0(mem_stage_inst_dmem_n210), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n370) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u343 ( .A(mem_stage_inst_dmem_n385), .B(
        mem_stage_inst_dmem_n375), .C(mem_stage_inst_dmem_n380), .D(
        mem_stage_inst_dmem_n370), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n390) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u342 ( .A(mem_stage_inst_dmem_n302), .B(
        mem_stage_inst_dmem_n303), .C(mem_stage_inst_dmem_n304), .D(
        mem_stage_inst_dmem_n305), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n301) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u341 ( .A(mem_stage_inst_dmem_n297), .B(
        mem_stage_inst_dmem_n298), .C(mem_stage_inst_dmem_n299), .D(
        mem_stage_inst_dmem_n300), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n296) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u340 ( .A(mem_stage_inst_dmem_n287), .B(
        mem_stage_inst_dmem_n288), .C(mem_stage_inst_dmem_n289), .D(
        mem_stage_inst_dmem_n290), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n286) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u339 ( .A(mem_stage_inst_dmem_n301), .B(
        mem_stage_inst_dmem_n291), .C(mem_stage_inst_dmem_n296), .D(
        mem_stage_inst_dmem_n286), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n306) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u338 ( .A(mem_stage_inst_dmem_n5618), 
        .B(mem_stage_inst_dmem_n5619), .C(mem_stage_inst_dmem_n5620), .D(
        mem_stage_inst_dmem_n5621), .S0(mem_stage_inst_dmem_n214), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5617) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u337 ( .A(mem_stage_inst_dmem_n5613), 
        .B(mem_stage_inst_dmem_n5614), .C(mem_stage_inst_dmem_n5615), .D(
        mem_stage_inst_dmem_n5616), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5612) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u336 ( .A(mem_stage_inst_dmem_n5603), 
        .B(mem_stage_inst_dmem_n5604), .C(mem_stage_inst_dmem_n5605), .D(
        mem_stage_inst_dmem_n5606), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5602) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u335 ( .A(mem_stage_inst_dmem_n5617), 
        .B(mem_stage_inst_dmem_n5607), .C(mem_stage_inst_dmem_n5612), .D(
        mem_stage_inst_dmem_n5602), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5663) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u334 ( .A(mem_stage_inst_dmem_n5534), 
        .B(mem_stage_inst_dmem_n5535), .C(mem_stage_inst_dmem_n5536), .D(
        mem_stage_inst_dmem_n5537), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5533) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u333 ( .A(mem_stage_inst_dmem_n5529), 
        .B(mem_stage_inst_dmem_n5530), .C(mem_stage_inst_dmem_n5531), .D(
        mem_stage_inst_dmem_n5532), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5528) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u332 ( .A(mem_stage_inst_dmem_n5519), 
        .B(mem_stage_inst_dmem_n5520), .C(mem_stage_inst_dmem_n5521), .D(
        mem_stage_inst_dmem_n5522), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5518) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u331 ( .A(mem_stage_inst_dmem_n5533), 
        .B(mem_stage_inst_dmem_n5523), .C(mem_stage_inst_dmem_n5528), .D(
        mem_stage_inst_dmem_n5518), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5579) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u330 ( .A(mem_stage_inst_dmem_n5450), 
        .B(mem_stage_inst_dmem_n5451), .C(mem_stage_inst_dmem_n5452), .D(
        mem_stage_inst_dmem_n5453), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n5449) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u329 ( .A(mem_stage_inst_dmem_n5445), 
        .B(mem_stage_inst_dmem_n5446), .C(mem_stage_inst_dmem_n5447), .D(
        mem_stage_inst_dmem_n5448), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5444) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u328 ( .A(mem_stage_inst_dmem_n5435), 
        .B(mem_stage_inst_dmem_n5436), .C(mem_stage_inst_dmem_n5437), .D(
        mem_stage_inst_dmem_n5438), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5434) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u327 ( .A(mem_stage_inst_dmem_n5449), 
        .B(mem_stage_inst_dmem_n5439), .C(mem_stage_inst_dmem_n5444), .D(
        mem_stage_inst_dmem_n5434), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5495) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u326 ( .A(mem_stage_inst_dmem_n5366), 
        .B(mem_stage_inst_dmem_n5367), .C(mem_stage_inst_dmem_n5368), .D(
        mem_stage_inst_dmem_n5369), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n5365) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u325 ( .A(mem_stage_inst_dmem_n5361), 
        .B(mem_stage_inst_dmem_n5362), .C(mem_stage_inst_dmem_n5363), .D(
        mem_stage_inst_dmem_n5364), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5360) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u324 ( .A(mem_stage_inst_dmem_n5351), 
        .B(mem_stage_inst_dmem_n5352), .C(mem_stage_inst_dmem_n5353), .D(
        mem_stage_inst_dmem_n5354), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5350) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u323 ( .A(mem_stage_inst_dmem_n5365), 
        .B(mem_stage_inst_dmem_n5355), .C(mem_stage_inst_dmem_n5360), .D(
        mem_stage_inst_dmem_n5350), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5411) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u322 ( .A(mem_stage_inst_dmem_n5282), 
        .B(mem_stage_inst_dmem_n5283), .C(mem_stage_inst_dmem_n5284), .D(
        mem_stage_inst_dmem_n5285), .S0(mem_stage_inst_dmem_n216), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5281) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u321 ( .A(mem_stage_inst_dmem_n5277), 
        .B(mem_stage_inst_dmem_n5278), .C(mem_stage_inst_dmem_n5279), .D(
        mem_stage_inst_dmem_n5280), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n5276) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u320 ( .A(mem_stage_inst_dmem_n5267), 
        .B(mem_stage_inst_dmem_n5268), .C(mem_stage_inst_dmem_n5269), .D(
        mem_stage_inst_dmem_n5270), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n5266) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u319 ( .A(mem_stage_inst_dmem_n5281), 
        .B(mem_stage_inst_dmem_n5271), .C(mem_stage_inst_dmem_n5276), .D(
        mem_stage_inst_dmem_n5266), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5327) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u318 ( .A(mem_stage_inst_dmem_n5198), 
        .B(mem_stage_inst_dmem_n5199), .C(mem_stage_inst_dmem_n5200), .D(
        mem_stage_inst_dmem_n5201), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5197) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u317 ( .A(mem_stage_inst_dmem_n5193), 
        .B(mem_stage_inst_dmem_n5194), .C(mem_stage_inst_dmem_n5195), .D(
        mem_stage_inst_dmem_n5196), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5192) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u316 ( .A(mem_stage_inst_dmem_n5183), 
        .B(mem_stage_inst_dmem_n5184), .C(mem_stage_inst_dmem_n5185), .D(
        mem_stage_inst_dmem_n5186), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5182) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u315 ( .A(mem_stage_inst_dmem_n5197), 
        .B(mem_stage_inst_dmem_n5187), .C(mem_stage_inst_dmem_n5192), .D(
        mem_stage_inst_dmem_n5182), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5243) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u314 ( .A(mem_stage_inst_dmem_n5114), 
        .B(mem_stage_inst_dmem_n5115), .C(mem_stage_inst_dmem_n5116), .D(
        mem_stage_inst_dmem_n5117), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5113) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u313 ( .A(mem_stage_inst_dmem_n5109), 
        .B(mem_stage_inst_dmem_n5110), .C(mem_stage_inst_dmem_n5111), .D(
        mem_stage_inst_dmem_n5112), .S0(mem_stage_inst_dmem_n214), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n5108) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u312 ( .A(mem_stage_inst_dmem_n5099), 
        .B(mem_stage_inst_dmem_n5100), .C(mem_stage_inst_dmem_n5101), .D(
        mem_stage_inst_dmem_n5102), .S0(mem_stage_inst_dmem_n214), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5098) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u311 ( .A(mem_stage_inst_dmem_n5113), 
        .B(mem_stage_inst_dmem_n5103), .C(mem_stage_inst_dmem_n5108), .D(
        mem_stage_inst_dmem_n5098), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5159) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u310 ( .A(mem_stage_inst_dmem_n5030), 
        .B(mem_stage_inst_dmem_n5031), .C(mem_stage_inst_dmem_n5032), .D(
        mem_stage_inst_dmem_n5033), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n5029) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u309 ( .A(mem_stage_inst_dmem_n5025), 
        .B(mem_stage_inst_dmem_n5026), .C(mem_stage_inst_dmem_n5027), .D(
        mem_stage_inst_dmem_n5028), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n5024) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u308 ( .A(mem_stage_inst_dmem_n5015), 
        .B(mem_stage_inst_dmem_n5016), .C(mem_stage_inst_dmem_n5017), .D(
        mem_stage_inst_dmem_n5018), .S0(mem_stage_inst_dmem_n213), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n5014) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u307 ( .A(mem_stage_inst_dmem_n5029), 
        .B(mem_stage_inst_dmem_n5019), .C(mem_stage_inst_dmem_n5024), .D(
        mem_stage_inst_dmem_n5014), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5075) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u306 ( .A(mem_stage_inst_dmem_n4946), 
        .B(mem_stage_inst_dmem_n4947), .C(mem_stage_inst_dmem_n4948), .D(
        mem_stage_inst_dmem_n4949), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4945) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u305 ( .A(mem_stage_inst_dmem_n4941), 
        .B(mem_stage_inst_dmem_n4942), .C(mem_stage_inst_dmem_n4943), .D(
        mem_stage_inst_dmem_n4944), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n4940) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u304 ( .A(mem_stage_inst_dmem_n4931), 
        .B(mem_stage_inst_dmem_n4932), .C(mem_stage_inst_dmem_n4933), .D(
        mem_stage_inst_dmem_n4934), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n4930) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u303 ( .A(mem_stage_inst_dmem_n4945), 
        .B(mem_stage_inst_dmem_n4935), .C(mem_stage_inst_dmem_n4940), .D(
        mem_stage_inst_dmem_n4930), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4991) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u302 ( .A(mem_stage_inst_dmem_n4862), 
        .B(mem_stage_inst_dmem_n4863), .C(mem_stage_inst_dmem_n4864), .D(
        mem_stage_inst_dmem_n4865), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4861) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u301 ( .A(mem_stage_inst_dmem_n4857), 
        .B(mem_stage_inst_dmem_n4858), .C(mem_stage_inst_dmem_n4859), .D(
        mem_stage_inst_dmem_n4860), .S0(ex_pipeline_reg_out[25]), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4856) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u300 ( .A(mem_stage_inst_dmem_n4847), 
        .B(mem_stage_inst_dmem_n4848), .C(mem_stage_inst_dmem_n4849), .D(
        mem_stage_inst_dmem_n4850), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n4846) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u299 ( .A(mem_stage_inst_dmem_n4861), 
        .B(mem_stage_inst_dmem_n4851), .C(mem_stage_inst_dmem_n4856), .D(
        mem_stage_inst_dmem_n4846), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4907) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u298 ( .A(mem_stage_inst_dmem_n4778), 
        .B(mem_stage_inst_dmem_n4779), .C(mem_stage_inst_dmem_n4780), .D(
        mem_stage_inst_dmem_n4781), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4777) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u297 ( .A(mem_stage_inst_dmem_n4773), 
        .B(mem_stage_inst_dmem_n4774), .C(mem_stage_inst_dmem_n4775), .D(
        mem_stage_inst_dmem_n4776), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4772) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u296 ( .A(mem_stage_inst_dmem_n4763), 
        .B(mem_stage_inst_dmem_n4764), .C(mem_stage_inst_dmem_n4765), .D(
        mem_stage_inst_dmem_n4766), .S0(mem_stage_inst_dmem_n215), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n4762) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u295 ( .A(mem_stage_inst_dmem_n4777), 
        .B(mem_stage_inst_dmem_n4767), .C(mem_stage_inst_dmem_n4772), .D(
        mem_stage_inst_dmem_n4762), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4823) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u294 ( .A(mem_stage_inst_dmem_n4694), 
        .B(mem_stage_inst_dmem_n4695), .C(mem_stage_inst_dmem_n4696), .D(
        mem_stage_inst_dmem_n4697), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4693) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u293 ( .A(mem_stage_inst_dmem_n4689), 
        .B(mem_stage_inst_dmem_n4690), .C(mem_stage_inst_dmem_n4691), .D(
        mem_stage_inst_dmem_n4692), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4688) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u292 ( .A(mem_stage_inst_dmem_n4679), 
        .B(mem_stage_inst_dmem_n4680), .C(mem_stage_inst_dmem_n4681), .D(
        mem_stage_inst_dmem_n4682), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n199), .Y(mem_stage_inst_dmem_n4678) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u291 ( .A(mem_stage_inst_dmem_n4693), 
        .B(mem_stage_inst_dmem_n4683), .C(mem_stage_inst_dmem_n4688), .D(
        mem_stage_inst_dmem_n4678), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4739) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u290 ( .A(mem_stage_inst_dmem_n514), .B(
        mem_stage_inst_dmem_n515), .C(mem_stage_inst_dmem_n516), .D(
        mem_stage_inst_dmem_n517), .S0(mem_stage_inst_dmem_n211), .S1(
        ex_pipeline_reg_out[24]), .Y(mem_stage_inst_dmem_n513) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u289 ( .A(mem_stage_inst_dmem_n509), .B(
        mem_stage_inst_dmem_n510), .C(mem_stage_inst_dmem_n511), .D(
        mem_stage_inst_dmem_n512), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n200), .Y(mem_stage_inst_dmem_n508) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u288 ( .A(mem_stage_inst_dmem_n499), .B(
        mem_stage_inst_dmem_n500), .C(mem_stage_inst_dmem_n501), .D(
        mem_stage_inst_dmem_n502), .S0(mem_stage_inst_dmem_n211), .S1(
        mem_stage_inst_dmem_n201), .Y(mem_stage_inst_dmem_n498) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u287 ( .A(mem_stage_inst_dmem_n513), .B(
        mem_stage_inst_dmem_n503), .C(mem_stage_inst_dmem_n508), .D(
        mem_stage_inst_dmem_n498), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n559) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u286 ( .A(mem_stage_inst_dmem_n430), .B(
        mem_stage_inst_dmem_n431), .C(mem_stage_inst_dmem_n432), .D(
        mem_stage_inst_dmem_n433), .S0(mem_stage_inst_dmem_n212), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n429) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u285 ( .A(mem_stage_inst_dmem_n425), .B(
        mem_stage_inst_dmem_n426), .C(mem_stage_inst_dmem_n427), .D(
        mem_stage_inst_dmem_n428), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n202), .Y(mem_stage_inst_dmem_n424) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u284 ( .A(mem_stage_inst_dmem_n415), .B(
        mem_stage_inst_dmem_n416), .C(mem_stage_inst_dmem_n417), .D(
        mem_stage_inst_dmem_n418), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n203), .Y(mem_stage_inst_dmem_n414) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u283 ( .A(mem_stage_inst_dmem_n429), .B(
        mem_stage_inst_dmem_n419), .C(mem_stage_inst_dmem_n424), .D(
        mem_stage_inst_dmem_n414), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n475) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u282 ( .A(mem_stage_inst_dmem_n346), .B(
        mem_stage_inst_dmem_n347), .C(mem_stage_inst_dmem_n348), .D(
        mem_stage_inst_dmem_n349), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n345) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u281 ( .A(mem_stage_inst_dmem_n341), .B(
        mem_stage_inst_dmem_n342), .C(mem_stage_inst_dmem_n343), .D(
        mem_stage_inst_dmem_n344), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n340) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u280 ( .A(mem_stage_inst_dmem_n331), .B(
        mem_stage_inst_dmem_n332), .C(mem_stage_inst_dmem_n333), .D(
        mem_stage_inst_dmem_n334), .S0(mem_stage_inst_dmem_n209), .S1(
        mem_stage_inst_dmem_n198), .Y(mem_stage_inst_dmem_n330) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u279 ( .A(mem_stage_inst_dmem_n345), .B(
        mem_stage_inst_dmem_n335), .C(mem_stage_inst_dmem_n340), .D(
        mem_stage_inst_dmem_n330), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n391) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u278 ( .A(mem_stage_inst_dmem_n262), .B(
        mem_stage_inst_dmem_n263), .C(mem_stage_inst_dmem_n264), .D(
        mem_stage_inst_dmem_n265), .S0(mem_stage_inst_dmem_n210), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n261) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u277 ( .A(mem_stage_inst_dmem_n257), .B(
        mem_stage_inst_dmem_n258), .C(mem_stage_inst_dmem_n259), .D(
        mem_stage_inst_dmem_n260), .S0(mem_stage_inst_dmem_n217), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n256) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u276 ( .A(mem_stage_inst_dmem_n247), .B(
        mem_stage_inst_dmem_n248), .C(mem_stage_inst_dmem_n249), .D(
        mem_stage_inst_dmem_n250), .S0(mem_stage_inst_dmem_n216), .S1(
        mem_stage_inst_dmem_n197), .Y(mem_stage_inst_dmem_n246) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u275 ( .A(mem_stage_inst_dmem_n261), .B(
        mem_stage_inst_dmem_n251), .C(mem_stage_inst_dmem_n256), .D(
        mem_stage_inst_dmem_n246), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n307) );
  INV_X1M_A12TS mem_stage_inst_dmem_u274 ( .A(ex_pipeline_reg_out[25]), .Y(
        mem_stage_inst_dmem_n225) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u273 ( .A(mem_stage_inst_dmem_n225), .Y(
        mem_stage_inst_dmem_n218) );
  INV_X1M_A12TS mem_stage_inst_dmem_u272 ( .A(ex_pipeline_reg_out[23]), .Y(
        mem_stage_inst_dmem_n196) );
  INV_X1M_A12TS mem_stage_inst_dmem_u271 ( .A(ex_pipeline_reg_out[22]), .Y(
        mem_stage_inst_dmem_n98) );
  INV_X1M_A12TS mem_stage_inst_dmem_u270 ( .A(ex_pipeline_reg_out[24]), .Y(
        mem_stage_inst_dmem_n208) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u269 ( .A(mem_stage_inst_dmem_n208), .Y(
        mem_stage_inst_dmem_n204) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u268 ( .A(mem_stage_inst_dmem_n5637), 
        .B(mem_stage_inst_dmem_n5627), .C(mem_stage_inst_dmem_n5632), .D(
        mem_stage_inst_dmem_n5622), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5664) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u267 ( .A(mem_stage_inst_dmem_n5597), 
        .B(mem_stage_inst_dmem_n5587), .C(mem_stage_inst_dmem_n5592), .D(
        mem_stage_inst_dmem_n5582), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5665) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u266 ( .A(mem_stage_inst_dmem_n5662), 
        .B(mem_stage_inst_dmem_n5663), .C(mem_stage_inst_dmem_n5664), .D(
        mem_stage_inst_dmem_n5665), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[15]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u265 ( .A(mem_stage_inst_dmem_n5553), 
        .B(mem_stage_inst_dmem_n5543), .C(mem_stage_inst_dmem_n5548), .D(
        mem_stage_inst_dmem_n5538), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5580) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u264 ( .A(mem_stage_inst_dmem_n5513), 
        .B(mem_stage_inst_dmem_n5503), .C(mem_stage_inst_dmem_n5508), .D(
        mem_stage_inst_dmem_n5498), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5581) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u263 ( .A(mem_stage_inst_dmem_n5578), 
        .B(mem_stage_inst_dmem_n5579), .C(mem_stage_inst_dmem_n5580), .D(
        mem_stage_inst_dmem_n5581), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[14]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u262 ( .A(mem_stage_inst_dmem_n5469), 
        .B(mem_stage_inst_dmem_n5459), .C(mem_stage_inst_dmem_n5464), .D(
        mem_stage_inst_dmem_n5454), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5496) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u261 ( .A(mem_stage_inst_dmem_n5429), 
        .B(mem_stage_inst_dmem_n5419), .C(mem_stage_inst_dmem_n5424), .D(
        mem_stage_inst_dmem_n5414), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5497) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u260 ( .A(mem_stage_inst_dmem_n5494), 
        .B(mem_stage_inst_dmem_n5495), .C(mem_stage_inst_dmem_n5496), .D(
        mem_stage_inst_dmem_n5497), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[13]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u259 ( .A(mem_stage_inst_dmem_n5385), 
        .B(mem_stage_inst_dmem_n5375), .C(mem_stage_inst_dmem_n5380), .D(
        mem_stage_inst_dmem_n5370), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5412) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u258 ( .A(mem_stage_inst_dmem_n5345), 
        .B(mem_stage_inst_dmem_n5335), .C(mem_stage_inst_dmem_n5340), .D(
        mem_stage_inst_dmem_n5330), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5413) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u257 ( .A(mem_stage_inst_dmem_n5410), 
        .B(mem_stage_inst_dmem_n5411), .C(mem_stage_inst_dmem_n5412), .D(
        mem_stage_inst_dmem_n5413), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[12]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u256 ( .A(mem_stage_inst_dmem_n5301), 
        .B(mem_stage_inst_dmem_n5291), .C(mem_stage_inst_dmem_n5296), .D(
        mem_stage_inst_dmem_n5286), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5328) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u255 ( .A(mem_stage_inst_dmem_n5261), 
        .B(mem_stage_inst_dmem_n5251), .C(mem_stage_inst_dmem_n5256), .D(
        mem_stage_inst_dmem_n5246), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5329) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u254 ( .A(mem_stage_inst_dmem_n5326), 
        .B(mem_stage_inst_dmem_n5327), .C(mem_stage_inst_dmem_n5328), .D(
        mem_stage_inst_dmem_n5329), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[11]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u253 ( .A(mem_stage_inst_dmem_n5217), 
        .B(mem_stage_inst_dmem_n5207), .C(mem_stage_inst_dmem_n5212), .D(
        mem_stage_inst_dmem_n5202), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5244) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u252 ( .A(mem_stage_inst_dmem_n5177), 
        .B(mem_stage_inst_dmem_n5167), .C(mem_stage_inst_dmem_n5172), .D(
        mem_stage_inst_dmem_n5162), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5245) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u251 ( .A(mem_stage_inst_dmem_n5242), 
        .B(mem_stage_inst_dmem_n5243), .C(mem_stage_inst_dmem_n5244), .D(
        mem_stage_inst_dmem_n5245), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[10]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u250 ( .A(mem_stage_inst_dmem_n5133), 
        .B(mem_stage_inst_dmem_n5123), .C(mem_stage_inst_dmem_n5128), .D(
        mem_stage_inst_dmem_n5118), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5160) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u249 ( .A(mem_stage_inst_dmem_n5093), 
        .B(mem_stage_inst_dmem_n5083), .C(mem_stage_inst_dmem_n5088), .D(
        mem_stage_inst_dmem_n5078), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5161) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u248 ( .A(mem_stage_inst_dmem_n5158), 
        .B(mem_stage_inst_dmem_n5159), .C(mem_stage_inst_dmem_n5160), .D(
        mem_stage_inst_dmem_n5161), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[9]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u247 ( .A(mem_stage_inst_dmem_n5049), 
        .B(mem_stage_inst_dmem_n5039), .C(mem_stage_inst_dmem_n5044), .D(
        mem_stage_inst_dmem_n5034), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5076) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u246 ( .A(mem_stage_inst_dmem_n5009), 
        .B(mem_stage_inst_dmem_n4999), .C(mem_stage_inst_dmem_n5004), .D(
        mem_stage_inst_dmem_n4994), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n5077) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u245 ( .A(mem_stage_inst_dmem_n5074), 
        .B(mem_stage_inst_dmem_n5075), .C(mem_stage_inst_dmem_n5076), .D(
        mem_stage_inst_dmem_n5077), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[8]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u244 ( .A(mem_stage_inst_dmem_n4965), 
        .B(mem_stage_inst_dmem_n4955), .C(mem_stage_inst_dmem_n4960), .D(
        mem_stage_inst_dmem_n4950), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4992) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u243 ( .A(mem_stage_inst_dmem_n4925), 
        .B(mem_stage_inst_dmem_n4915), .C(mem_stage_inst_dmem_n4920), .D(
        mem_stage_inst_dmem_n4910), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4993) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u242 ( .A(mem_stage_inst_dmem_n4990), 
        .B(mem_stage_inst_dmem_n4991), .C(mem_stage_inst_dmem_n4992), .D(
        mem_stage_inst_dmem_n4993), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[7]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u241 ( .A(mem_stage_inst_dmem_n4881), 
        .B(mem_stage_inst_dmem_n4871), .C(mem_stage_inst_dmem_n4876), .D(
        mem_stage_inst_dmem_n4866), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4908) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u240 ( .A(mem_stage_inst_dmem_n4841), 
        .B(mem_stage_inst_dmem_n4831), .C(mem_stage_inst_dmem_n4836), .D(
        mem_stage_inst_dmem_n4826), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4909) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u239 ( .A(mem_stage_inst_dmem_n4906), 
        .B(mem_stage_inst_dmem_n4907), .C(mem_stage_inst_dmem_n4908), .D(
        mem_stage_inst_dmem_n4909), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[6]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u238 ( .A(mem_stage_inst_dmem_n4797), 
        .B(mem_stage_inst_dmem_n4787), .C(mem_stage_inst_dmem_n4792), .D(
        mem_stage_inst_dmem_n4782), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4824) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u237 ( .A(mem_stage_inst_dmem_n4757), 
        .B(mem_stage_inst_dmem_n4747), .C(mem_stage_inst_dmem_n4752), .D(
        mem_stage_inst_dmem_n4742), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4825) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u236 ( .A(mem_stage_inst_dmem_n4822), 
        .B(mem_stage_inst_dmem_n4823), .C(mem_stage_inst_dmem_n4824), .D(
        mem_stage_inst_dmem_n4825), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[5]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u235 ( .A(mem_stage_inst_dmem_n4713), 
        .B(mem_stage_inst_dmem_n4703), .C(mem_stage_inst_dmem_n4708), .D(
        mem_stage_inst_dmem_n4698), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4740) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u234 ( .A(mem_stage_inst_dmem_n4673), 
        .B(mem_stage_inst_dmem_n4663), .C(mem_stage_inst_dmem_n4668), .D(
        mem_stage_inst_dmem_n562), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n4741) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u233 ( .A(mem_stage_inst_dmem_n4738), 
        .B(mem_stage_inst_dmem_n4739), .C(mem_stage_inst_dmem_n4740), .D(
        mem_stage_inst_dmem_n4741), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[4]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u232 ( .A(mem_stage_inst_dmem_n533), .B(
        mem_stage_inst_dmem_n523), .C(mem_stage_inst_dmem_n528), .D(
        mem_stage_inst_dmem_n518), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n560) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u231 ( .A(mem_stage_inst_dmem_n493), .B(
        mem_stage_inst_dmem_n483), .C(mem_stage_inst_dmem_n488), .D(
        mem_stage_inst_dmem_n478), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n561) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u230 ( .A(mem_stage_inst_dmem_n558), .B(
        mem_stage_inst_dmem_n559), .C(mem_stage_inst_dmem_n560), .D(
        mem_stage_inst_dmem_n561), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[3]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u229 ( .A(mem_stage_inst_dmem_n449), .B(
        mem_stage_inst_dmem_n439), .C(mem_stage_inst_dmem_n444), .D(
        mem_stage_inst_dmem_n434), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n476) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u228 ( .A(mem_stage_inst_dmem_n409), .B(
        mem_stage_inst_dmem_n399), .C(mem_stage_inst_dmem_n404), .D(
        mem_stage_inst_dmem_n394), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n477) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u227 ( .A(mem_stage_inst_dmem_n474), .B(
        mem_stage_inst_dmem_n475), .C(mem_stage_inst_dmem_n476), .D(
        mem_stage_inst_dmem_n477), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[2]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u226 ( .A(mem_stage_inst_dmem_n365), .B(
        mem_stage_inst_dmem_n355), .C(mem_stage_inst_dmem_n360), .D(
        mem_stage_inst_dmem_n350), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n392) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u225 ( .A(mem_stage_inst_dmem_n325), .B(
        mem_stage_inst_dmem_n315), .C(mem_stage_inst_dmem_n320), .D(
        mem_stage_inst_dmem_n310), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n393) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u224 ( .A(mem_stage_inst_dmem_n390), .B(
        mem_stage_inst_dmem_n391), .C(mem_stage_inst_dmem_n392), .D(
        mem_stage_inst_dmem_n393), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[1]) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u223 ( .A(mem_stage_inst_dmem_n281), .B(
        mem_stage_inst_dmem_n271), .C(mem_stage_inst_dmem_n276), .D(
        mem_stage_inst_dmem_n266), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n308) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u222 ( .A(mem_stage_inst_dmem_n241), .B(
        mem_stage_inst_dmem_n231), .C(mem_stage_inst_dmem_n236), .D(
        mem_stage_inst_dmem_n226), .S0(ex_pipeline_reg_out[27]), .S1(
        ex_pipeline_reg_out[26]), .Y(mem_stage_inst_dmem_n309) );
  MXIT4_X1M_A12TS mem_stage_inst_dmem_u221 ( .A(mem_stage_inst_dmem_n306), .B(
        mem_stage_inst_dmem_n307), .C(mem_stage_inst_dmem_n308), .D(
        mem_stage_inst_dmem_n309), .S0(ex_pipeline_reg_out[29]), .S1(
        ex_pipeline_reg_out[28]), .Y(mem_stage_inst_mem_read_data[0]) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u220 ( .A(mem_stage_inst_dmem_n98), .Y(
        mem_stage_inst_dmem_n95) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u219 ( .A(mem_stage_inst_dmem_n96), .Y(
        mem_stage_inst_dmem_n94) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u218 ( .A(mem_stage_inst_dmem_n196), .Y(
        mem_stage_inst_dmem_n190) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u217 ( .A(mem_stage_inst_dmem_n196), .Y(
        mem_stage_inst_dmem_n191) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u216 ( .A(mem_stage_inst_dmem_n89), .Y(
        mem_stage_inst_dmem_n93) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u215 ( .A(mem_stage_inst_dmem_n88), .Y(
        mem_stage_inst_dmem_n97) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u214 ( .A(mem_stage_inst_dmem_n194), .Y(
        mem_stage_inst_dmem_n188) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u213 ( .A(mem_stage_inst_dmem_n88), .Y(
        mem_stage_inst_dmem_n96) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u212 ( .A(mem_stage_inst_dmem_n193), .Y(
        mem_stage_inst_dmem_n189) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u211 ( .A(mem_stage_inst_dmem_n98), .Y(
        mem_stage_inst_dmem_n90) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u210 ( .A(mem_stage_inst_dmem_n192), .Y(
        mem_stage_inst_dmem_n194) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u209 ( .A(mem_stage_inst_dmem_n98), .Y(
        mem_stage_inst_dmem_n91) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u208 ( .A(mem_stage_inst_dmem_n196), .Y(
        mem_stage_inst_dmem_n193) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u207 ( .A(mem_stage_inst_dmem_n98), .Y(
        mem_stage_inst_dmem_n89) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u206 ( .A(mem_stage_inst_dmem_n187), .Y(
        mem_stage_inst_dmem_n195) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u205 ( .A(mem_stage_inst_dmem_n95), .Y(
        mem_stage_inst_dmem_n92) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u204 ( .A(mem_stage_inst_dmem_n196), .Y(
        mem_stage_inst_dmem_n192) );
  INV_X1M_A12TS mem_stage_inst_dmem_u203 ( .A(mem_stage_inst_dmem_n204), .Y(
        mem_stage_inst_dmem_n198) );
  INV_X1M_A12TS mem_stage_inst_dmem_u202 ( .A(mem_stage_inst_dmem_n204), .Y(
        mem_stage_inst_dmem_n197) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u201 ( .A(mem_stage_inst_dmem_n225), .Y(
        mem_stage_inst_dmem_n219) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u200 ( .A(mem_stage_inst_dmem_n225), .Y(
        mem_stage_inst_dmem_n220) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u199 ( .A(mem_stage_inst_dmem_n222), .Y(
        mem_stage_inst_dmem_n221) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u198 ( .A(mem_stage_inst_dmem_n208), .Y(
        mem_stage_inst_dmem_n207) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u197 ( .A(mem_stage_inst_dmem_n208), .Y(
        mem_stage_inst_dmem_n206) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u196 ( .A(mem_stage_inst_dmem_n207), .Y(
        mem_stage_inst_dmem_n205) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u195 ( .A(mem_stage_inst_dmem_n225), .Y(
        mem_stage_inst_dmem_n222) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u194 ( .A(mem_stage_inst_dmem_n219), .Y(
        mem_stage_inst_dmem_n223) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u193 ( .A(mem_stage_inst_dmem_n220), .Y(
        mem_stage_inst_dmem_n224) );
  INV_X1M_A12TS mem_stage_inst_dmem_u192 ( .A(mem_stage_inst_dmem_n207), .Y(
        mem_stage_inst_dmem_n203) );
  INV_X1M_A12TS mem_stage_inst_dmem_u191 ( .A(mem_stage_inst_dmem_n207), .Y(
        mem_stage_inst_dmem_n202) );
  INV_X1M_A12TS mem_stage_inst_dmem_u190 ( .A(mem_stage_inst_dmem_n206), .Y(
        mem_stage_inst_dmem_n201) );
  INV_X1M_A12TS mem_stage_inst_dmem_u189 ( .A(mem_stage_inst_dmem_n206), .Y(
        mem_stage_inst_dmem_n200) );
  INV_X1M_A12TS mem_stage_inst_dmem_u188 ( .A(mem_stage_inst_dmem_n205), .Y(
        mem_stage_inst_dmem_n199) );
  INV_X1M_A12TS mem_stage_inst_dmem_u187 ( .A(mem_stage_inst_dmem_n219), .Y(
        mem_stage_inst_dmem_n216) );
  INV_X1M_A12TS mem_stage_inst_dmem_u186 ( .A(mem_stage_inst_dmem_n219), .Y(
        mem_stage_inst_dmem_n217) );
  INV_X1M_A12TS mem_stage_inst_dmem_u185 ( .A(mem_stage_inst_dmem_n220), .Y(
        mem_stage_inst_dmem_n215) );
  INV_X1M_A12TS mem_stage_inst_dmem_u184 ( .A(mem_stage_inst_dmem_n221), .Y(
        mem_stage_inst_dmem_n214) );
  INV_X1M_A12TS mem_stage_inst_dmem_u183 ( .A(mem_stage_inst_dmem_n221), .Y(
        mem_stage_inst_dmem_n213) );
  INV_X1M_A12TS mem_stage_inst_dmem_u182 ( .A(mem_stage_inst_dmem_n222), .Y(
        mem_stage_inst_dmem_n211) );
  INV_X1M_A12TS mem_stage_inst_dmem_u181 ( .A(mem_stage_inst_dmem_n222), .Y(
        mem_stage_inst_dmem_n212) );
  INV_X1M_A12TS mem_stage_inst_dmem_u180 ( .A(mem_stage_inst_dmem_n223), .Y(
        mem_stage_inst_dmem_n210) );
  INV_X1M_A12TS mem_stage_inst_dmem_u179 ( .A(mem_stage_inst_dmem_n224), .Y(
        mem_stage_inst_dmem_n209) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u178 ( .A(mem_stage_inst_dmem_n188), .Y(
        mem_stage_inst_dmem_n187) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u177 ( .A(mem_stage_inst_dmem_n89), .Y(
        mem_stage_inst_dmem_n88) );
  INV_X1M_A12TS mem_stage_inst_dmem_u176 ( .A(mem_stage_inst_dmem_n88), .Y(
        mem_stage_inst_dmem_n64) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u175 ( .A(mem_stage_inst_dmem_n190), .Y(
        mem_stage_inst_dmem_n181) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u174 ( .A(mem_stage_inst_dmem_n95), .Y(
        mem_stage_inst_dmem_n72) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u173 ( .A(mem_stage_inst_dmem_n190), .Y(
        mem_stage_inst_dmem_n180) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u172 ( .A(mem_stage_inst_dmem_n191), .Y(
        mem_stage_inst_dmem_n179) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u171 ( .A(mem_stage_inst_dmem_n93), .Y(
        mem_stage_inst_dmem_n74) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u170 ( .A(mem_stage_inst_dmem_n191), .Y(
        mem_stage_inst_dmem_n178) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u169 ( .A(mem_stage_inst_dmem_n93), .Y(
        mem_stage_inst_dmem_n75) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u168 ( .A(mem_stage_inst_dmem_n94), .Y(
        mem_stage_inst_dmem_n73) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u167 ( .A(mem_stage_inst_dmem_n188), .Y(
        mem_stage_inst_dmem_n185) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u166 ( .A(mem_stage_inst_dmem_n189), .Y(
        mem_stage_inst_dmem_n184) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u165 ( .A(mem_stage_inst_dmem_n188), .Y(
        mem_stage_inst_dmem_n186) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u164 ( .A(mem_stage_inst_dmem_n96), .Y(
        mem_stage_inst_dmem_n71) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u163 ( .A(mem_stage_inst_dmem_n189), .Y(
        mem_stage_inst_dmem_n182) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u162 ( .A(mem_stage_inst_dmem_n189), .Y(
        mem_stage_inst_dmem_n183) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u161 ( .A(mem_stage_inst_dmem_n90), .Y(
        mem_stage_inst_dmem_n84) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u160 ( .A(mem_stage_inst_dmem_n90), .Y(
        mem_stage_inst_dmem_n85) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u159 ( .A(mem_stage_inst_dmem_n91), .Y(
        mem_stage_inst_dmem_n82) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u158 ( .A(mem_stage_inst_dmem_n90), .Y(
        mem_stage_inst_dmem_n83) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u157 ( .A(mem_stage_inst_dmem_n89), .Y(
        mem_stage_inst_dmem_n87) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u156 ( .A(mem_stage_inst_dmem_n92), .Y(
        mem_stage_inst_dmem_n78) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u155 ( .A(mem_stage_inst_dmem_n192), .Y(
        mem_stage_inst_dmem_n175) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u154 ( .A(mem_stage_inst_dmem_n89), .Y(
        mem_stage_inst_dmem_n86) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u153 ( .A(mem_stage_inst_dmem_n92), .Y(
        mem_stage_inst_dmem_n77) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u152 ( .A(mem_stage_inst_dmem_n192), .Y(
        mem_stage_inst_dmem_n176) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u151 ( .A(mem_stage_inst_dmem_n93), .Y(
        mem_stage_inst_dmem_n76) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u150 ( .A(mem_stage_inst_dmem_n191), .Y(
        mem_stage_inst_dmem_n177) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u149 ( .A(mem_stage_inst_dmem_n91), .Y(
        mem_stage_inst_dmem_n80) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u148 ( .A(mem_stage_inst_dmem_n193), .Y(
        mem_stage_inst_dmem_n173) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u147 ( .A(mem_stage_inst_dmem_n91), .Y(
        mem_stage_inst_dmem_n81) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u146 ( .A(mem_stage_inst_dmem_n92), .Y(
        mem_stage_inst_dmem_n79) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u145 ( .A(mem_stage_inst_dmem_n192), .Y(
        mem_stage_inst_dmem_n174) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u144 ( .A(mem_stage_inst_dmem_n96), .Y(
        mem_stage_inst_dmem_n69) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u143 ( .A(mem_stage_inst_dmem_n96), .Y(
        mem_stage_inst_dmem_n70) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u142 ( .A(mem_stage_inst_dmem_n193), .Y(
        mem_stage_inst_dmem_n171) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u141 ( .A(mem_stage_inst_dmem_n193), .Y(
        mem_stage_inst_dmem_n172) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u140 ( .A(mem_stage_inst_dmem_n195), .Y(
        mem_stage_inst_dmem_n165) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u139 ( .A(mem_stage_inst_dmem_n97), .Y(
        mem_stage_inst_dmem_n68) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u138 ( .A(mem_stage_inst_dmem_n97), .Y(
        mem_stage_inst_dmem_n67) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u137 ( .A(mem_stage_inst_dmem_n194), .Y(
        mem_stage_inst_dmem_n170) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u136 ( .A(mem_stage_inst_dmem_n194), .Y(
        mem_stage_inst_dmem_n169) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u135 ( .A(mem_stage_inst_dmem_n194), .Y(
        mem_stage_inst_dmem_n168) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u134 ( .A(mem_stage_inst_dmem_n195), .Y(
        mem_stage_inst_dmem_n167) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u133 ( .A(mem_stage_inst_dmem_n195), .Y(
        mem_stage_inst_dmem_n166) );
  BUFH_X1M_A12TS mem_stage_inst_dmem_u132 ( .A(mem_stage_inst_dmem_n97), .Y(
        mem_stage_inst_dmem_n66) );
  INV_X1M_A12TS mem_stage_inst_dmem_u131 ( .A(mem_stage_inst_dmem_n72), .Y(
        mem_stage_inst_dmem_n20) );
  INV_X1M_A12TS mem_stage_inst_dmem_u130 ( .A(mem_stage_inst_dmem_n72), .Y(
        mem_stage_inst_dmem_n21) );
  INV_X1M_A12TS mem_stage_inst_dmem_u129 ( .A(mem_stage_inst_dmem_n72), .Y(
        mem_stage_inst_dmem_n19) );
  INV_X1M_A12TS mem_stage_inst_dmem_u128 ( .A(mem_stage_inst_dmem_n74), .Y(
        mem_stage_inst_dmem_n25) );
  INV_X1M_A12TS mem_stage_inst_dmem_u127 ( .A(mem_stage_inst_dmem_n74), .Y(
        mem_stage_inst_dmem_n26) );
  INV_X1M_A12TS mem_stage_inst_dmem_u126 ( .A(mem_stage_inst_dmem_n75), .Y(
        mem_stage_inst_dmem_n27) );
  INV_X1M_A12TS mem_stage_inst_dmem_u125 ( .A(mem_stage_inst_dmem_n73), .Y(
        mem_stage_inst_dmem_n22) );
  INV_X1M_A12TS mem_stage_inst_dmem_u124 ( .A(mem_stage_inst_dmem_n73), .Y(
        mem_stage_inst_dmem_n23) );
  INV_X1M_A12TS mem_stage_inst_dmem_u123 ( .A(mem_stage_inst_dmem_n73), .Y(
        mem_stage_inst_dmem_n24) );
  INV_X1M_A12TS mem_stage_inst_dmem_u122 ( .A(mem_stage_inst_dmem_n71), .Y(
        mem_stage_inst_dmem_n15) );
  INV_X1M_A12TS mem_stage_inst_dmem_u121 ( .A(mem_stage_inst_dmem_n75), .Y(
        mem_stage_inst_dmem_n16) );
  INV_X1M_A12TS mem_stage_inst_dmem_u120 ( .A(mem_stage_inst_dmem_n71), .Y(
        mem_stage_inst_dmem_n18) );
  INV_X1M_A12TS mem_stage_inst_dmem_u119 ( .A(mem_stage_inst_dmem_n71), .Y(
        mem_stage_inst_dmem_n17) );
  INV_X1M_A12TS mem_stage_inst_dmem_u118 ( .A(mem_stage_inst_dmem_n84), .Y(
        mem_stage_inst_dmem_n52) );
  INV_X1M_A12TS mem_stage_inst_dmem_u117 ( .A(mem_stage_inst_dmem_n84), .Y(
        mem_stage_inst_dmem_n53) );
  INV_X1M_A12TS mem_stage_inst_dmem_u116 ( .A(mem_stage_inst_dmem_n84), .Y(
        mem_stage_inst_dmem_n54) );
  INV_X1M_A12TS mem_stage_inst_dmem_u115 ( .A(mem_stage_inst_dmem_n85), .Y(
        mem_stage_inst_dmem_n55) );
  INV_X1M_A12TS mem_stage_inst_dmem_u114 ( .A(mem_stage_inst_dmem_n85), .Y(
        mem_stage_inst_dmem_n56) );
  INV_X1M_A12TS mem_stage_inst_dmem_u113 ( .A(mem_stage_inst_dmem_n82), .Y(
        mem_stage_inst_dmem_n47) );
  INV_X1M_A12TS mem_stage_inst_dmem_u112 ( .A(mem_stage_inst_dmem_n82), .Y(
        mem_stage_inst_dmem_n48) );
  INV_X1M_A12TS mem_stage_inst_dmem_u111 ( .A(mem_stage_inst_dmem_n82), .Y(
        mem_stage_inst_dmem_n49) );
  INV_X1M_A12TS mem_stage_inst_dmem_u110 ( .A(mem_stage_inst_dmem_n83), .Y(
        mem_stage_inst_dmem_n50) );
  INV_X1M_A12TS mem_stage_inst_dmem_u109 ( .A(mem_stage_inst_dmem_n83), .Y(
        mem_stage_inst_dmem_n51) );
  INV_X1M_A12TS mem_stage_inst_dmem_u108 ( .A(mem_stage_inst_dmem_n87), .Y(
        mem_stage_inst_dmem_n61) );
  INV_X1M_A12TS mem_stage_inst_dmem_u107 ( .A(mem_stage_inst_dmem_n87), .Y(
        mem_stage_inst_dmem_n62) );
  INV_X1M_A12TS mem_stage_inst_dmem_u106 ( .A(mem_stage_inst_dmem_n87), .Y(
        mem_stage_inst_dmem_n63) );
  INV_X1M_A12TS mem_stage_inst_dmem_u105 ( .A(mem_stage_inst_dmem_n83), .Y(
        mem_stage_inst_dmem_n65) );
  INV_X1M_A12TS mem_stage_inst_dmem_u104 ( .A(mem_stage_inst_dmem_n78), .Y(
        mem_stage_inst_dmem_n37) );
  INV_X1M_A12TS mem_stage_inst_dmem_u103 ( .A(mem_stage_inst_dmem_n85), .Y(
        mem_stage_inst_dmem_n57) );
  INV_X1M_A12TS mem_stage_inst_dmem_u102 ( .A(mem_stage_inst_dmem_n86), .Y(
        mem_stage_inst_dmem_n58) );
  INV_X1M_A12TS mem_stage_inst_dmem_u101 ( .A(mem_stage_inst_dmem_n86), .Y(
        mem_stage_inst_dmem_n59) );
  INV_X1M_A12TS mem_stage_inst_dmem_u100 ( .A(mem_stage_inst_dmem_n86), .Y(
        mem_stage_inst_dmem_n60) );
  INV_X1M_A12TS mem_stage_inst_dmem_u99 ( .A(mem_stage_inst_dmem_n77), .Y(
        mem_stage_inst_dmem_n32) );
  INV_X1M_A12TS mem_stage_inst_dmem_u98 ( .A(mem_stage_inst_dmem_n77), .Y(
        mem_stage_inst_dmem_n33) );
  INV_X1M_A12TS mem_stage_inst_dmem_u97 ( .A(mem_stage_inst_dmem_n77), .Y(
        mem_stage_inst_dmem_n34) );
  INV_X1M_A12TS mem_stage_inst_dmem_u96 ( .A(mem_stage_inst_dmem_n78), .Y(
        mem_stage_inst_dmem_n35) );
  INV_X1M_A12TS mem_stage_inst_dmem_u95 ( .A(mem_stage_inst_dmem_n78), .Y(
        mem_stage_inst_dmem_n36) );
  INV_X1M_A12TS mem_stage_inst_dmem_u94 ( .A(mem_stage_inst_dmem_n75), .Y(
        mem_stage_inst_dmem_n28) );
  INV_X1M_A12TS mem_stage_inst_dmem_u93 ( .A(mem_stage_inst_dmem_n76), .Y(
        mem_stage_inst_dmem_n29) );
  INV_X1M_A12TS mem_stage_inst_dmem_u92 ( .A(mem_stage_inst_dmem_n76), .Y(
        mem_stage_inst_dmem_n30) );
  INV_X1M_A12TS mem_stage_inst_dmem_u91 ( .A(mem_stage_inst_dmem_n76), .Y(
        mem_stage_inst_dmem_n31) );
  INV_X1M_A12TS mem_stage_inst_dmem_u90 ( .A(mem_stage_inst_dmem_n80), .Y(
        mem_stage_inst_dmem_n42) );
  INV_X1M_A12TS mem_stage_inst_dmem_u89 ( .A(mem_stage_inst_dmem_n80), .Y(
        mem_stage_inst_dmem_n43) );
  INV_X1M_A12TS mem_stage_inst_dmem_u88 ( .A(mem_stage_inst_dmem_n81), .Y(
        mem_stage_inst_dmem_n44) );
  INV_X1M_A12TS mem_stage_inst_dmem_u87 ( .A(mem_stage_inst_dmem_n81), .Y(
        mem_stage_inst_dmem_n45) );
  INV_X1M_A12TS mem_stage_inst_dmem_u86 ( .A(mem_stage_inst_dmem_n81), .Y(
        mem_stage_inst_dmem_n46) );
  INV_X1M_A12TS mem_stage_inst_dmem_u85 ( .A(mem_stage_inst_dmem_n79), .Y(
        mem_stage_inst_dmem_n38) );
  INV_X1M_A12TS mem_stage_inst_dmem_u84 ( .A(mem_stage_inst_dmem_n79), .Y(
        mem_stage_inst_dmem_n39) );
  INV_X1M_A12TS mem_stage_inst_dmem_u83 ( .A(mem_stage_inst_dmem_n79), .Y(
        mem_stage_inst_dmem_n40) );
  INV_X1M_A12TS mem_stage_inst_dmem_u82 ( .A(mem_stage_inst_dmem_n80), .Y(
        mem_stage_inst_dmem_n41) );
  INV_X1M_A12TS mem_stage_inst_dmem_u81 ( .A(mem_stage_inst_dmem_n68), .Y(
        mem_stage_inst_dmem_n6) );
  INV_X1M_A12TS mem_stage_inst_dmem_u80 ( .A(mem_stage_inst_dmem_n68), .Y(
        mem_stage_inst_dmem_n7) );
  INV_X1M_A12TS mem_stage_inst_dmem_u79 ( .A(mem_stage_inst_dmem_n68), .Y(
        mem_stage_inst_dmem_n8) );
  INV_X1M_A12TS mem_stage_inst_dmem_u78 ( .A(mem_stage_inst_dmem_n69), .Y(
        mem_stage_inst_dmem_n9) );
  INV_X1M_A12TS mem_stage_inst_dmem_u77 ( .A(mem_stage_inst_dmem_n69), .Y(
        mem_stage_inst_dmem_n10) );
  INV_X1M_A12TS mem_stage_inst_dmem_u76 ( .A(mem_stage_inst_dmem_n67), .Y(
        mem_stage_inst_dmem_n5) );
  INV_X1M_A12TS mem_stage_inst_dmem_u75 ( .A(mem_stage_inst_dmem_n67), .Y(
        mem_stage_inst_dmem_n3) );
  INV_X1M_A12TS mem_stage_inst_dmem_u74 ( .A(mem_stage_inst_dmem_n67), .Y(
        mem_stage_inst_dmem_n4) );
  INV_X1M_A12TS mem_stage_inst_dmem_u73 ( .A(mem_stage_inst_dmem_n69), .Y(
        mem_stage_inst_dmem_n11) );
  INV_X1M_A12TS mem_stage_inst_dmem_u72 ( .A(mem_stage_inst_dmem_n70), .Y(
        mem_stage_inst_dmem_n13) );
  INV_X1M_A12TS mem_stage_inst_dmem_u71 ( .A(mem_stage_inst_dmem_n70), .Y(
        mem_stage_inst_dmem_n14) );
  INV_X1M_A12TS mem_stage_inst_dmem_u70 ( .A(mem_stage_inst_dmem_n70), .Y(
        mem_stage_inst_dmem_n12) );
  INV_X1M_A12TS mem_stage_inst_dmem_u69 ( .A(mem_stage_inst_dmem_n66), .Y(
        mem_stage_inst_dmem_n1) );
  INV_X1M_A12TS mem_stage_inst_dmem_u68 ( .A(mem_stage_inst_dmem_n66), .Y(
        mem_stage_inst_dmem_n2) );
  INV_X1M_A12TS mem_stage_inst_dmem_u67 ( .A(mem_stage_inst_dmem_n187), .Y(
        mem_stage_inst_dmem_n99) );
  INV_X1M_A12TS mem_stage_inst_dmem_u66 ( .A(mem_stage_inst_dmem_n187), .Y(
        mem_stage_inst_dmem_n100) );
  INV_X1M_A12TS mem_stage_inst_dmem_u65 ( .A(mem_stage_inst_dmem_n165), .Y(
        mem_stage_inst_dmem_n164) );
  INV_X1M_A12TS mem_stage_inst_dmem_u64 ( .A(mem_stage_inst_dmem_n181), .Y(
        mem_stage_inst_dmem_n116) );
  INV_X1M_A12TS mem_stage_inst_dmem_u63 ( .A(mem_stage_inst_dmem_n179), .Y(
        mem_stage_inst_dmem_n121) );
  INV_X1M_A12TS mem_stage_inst_dmem_u62 ( .A(mem_stage_inst_dmem_n179), .Y(
        mem_stage_inst_dmem_n122) );
  INV_X1M_A12TS mem_stage_inst_dmem_u61 ( .A(mem_stage_inst_dmem_n179), .Y(
        mem_stage_inst_dmem_n123) );
  INV_X1M_A12TS mem_stage_inst_dmem_u60 ( .A(mem_stage_inst_dmem_n178), .Y(
        mem_stage_inst_dmem_n124) );
  INV_X1M_A12TS mem_stage_inst_dmem_u59 ( .A(mem_stage_inst_dmem_n178), .Y(
        mem_stage_inst_dmem_n125) );
  INV_X1M_A12TS mem_stage_inst_dmem_u58 ( .A(mem_stage_inst_dmem_n181), .Y(
        mem_stage_inst_dmem_n117) );
  INV_X1M_A12TS mem_stage_inst_dmem_u57 ( .A(mem_stage_inst_dmem_n181), .Y(
        mem_stage_inst_dmem_n118) );
  INV_X1M_A12TS mem_stage_inst_dmem_u56 ( .A(mem_stage_inst_dmem_n180), .Y(
        mem_stage_inst_dmem_n119) );
  INV_X1M_A12TS mem_stage_inst_dmem_u55 ( .A(mem_stage_inst_dmem_n180), .Y(
        mem_stage_inst_dmem_n120) );
  INV_X1M_A12TS mem_stage_inst_dmem_u54 ( .A(mem_stage_inst_dmem_n185), .Y(
        mem_stage_inst_dmem_n104) );
  INV_X1M_A12TS mem_stage_inst_dmem_u53 ( .A(mem_stage_inst_dmem_n185), .Y(
        mem_stage_inst_dmem_n105) );
  INV_X1M_A12TS mem_stage_inst_dmem_u52 ( .A(mem_stage_inst_dmem_n185), .Y(
        mem_stage_inst_dmem_n106) );
  INV_X1M_A12TS mem_stage_inst_dmem_u51 ( .A(mem_stage_inst_dmem_n184), .Y(
        mem_stage_inst_dmem_n107) );
  INV_X1M_A12TS mem_stage_inst_dmem_u50 ( .A(mem_stage_inst_dmem_n184), .Y(
        mem_stage_inst_dmem_n108) );
  INV_X1M_A12TS mem_stage_inst_dmem_u49 ( .A(mem_stage_inst_dmem_n186), .Y(
        mem_stage_inst_dmem_n103) );
  INV_X1M_A12TS mem_stage_inst_dmem_u48 ( .A(mem_stage_inst_dmem_n186), .Y(
        mem_stage_inst_dmem_n101) );
  INV_X1M_A12TS mem_stage_inst_dmem_u47 ( .A(mem_stage_inst_dmem_n186), .Y(
        mem_stage_inst_dmem_n102) );
  INV_X1M_A12TS mem_stage_inst_dmem_u46 ( .A(mem_stage_inst_dmem_n182), .Y(
        mem_stage_inst_dmem_n113) );
  INV_X1M_A12TS mem_stage_inst_dmem_u45 ( .A(mem_stage_inst_dmem_n182), .Y(
        mem_stage_inst_dmem_n114) );
  INV_X1M_A12TS mem_stage_inst_dmem_u44 ( .A(mem_stage_inst_dmem_n182), .Y(
        mem_stage_inst_dmem_n115) );
  INV_X1M_A12TS mem_stage_inst_dmem_u43 ( .A(mem_stage_inst_dmem_n184), .Y(
        mem_stage_inst_dmem_n109) );
  INV_X1M_A12TS mem_stage_inst_dmem_u42 ( .A(mem_stage_inst_dmem_n183), .Y(
        mem_stage_inst_dmem_n111) );
  INV_X1M_A12TS mem_stage_inst_dmem_u41 ( .A(mem_stage_inst_dmem_n183), .Y(
        mem_stage_inst_dmem_n112) );
  INV_X1M_A12TS mem_stage_inst_dmem_u40 ( .A(mem_stage_inst_dmem_n183), .Y(
        mem_stage_inst_dmem_n110) );
  INV_X1M_A12TS mem_stage_inst_dmem_u39 ( .A(mem_stage_inst_dmem_n175), .Y(
        mem_stage_inst_dmem_n135) );
  INV_X1M_A12TS mem_stage_inst_dmem_u38 ( .A(mem_stage_inst_dmem_n176), .Y(
        mem_stage_inst_dmem_n130) );
  INV_X1M_A12TS mem_stage_inst_dmem_u37 ( .A(mem_stage_inst_dmem_n176), .Y(
        mem_stage_inst_dmem_n131) );
  INV_X1M_A12TS mem_stage_inst_dmem_u36 ( .A(mem_stage_inst_dmem_n176), .Y(
        mem_stage_inst_dmem_n132) );
  INV_X1M_A12TS mem_stage_inst_dmem_u35 ( .A(mem_stage_inst_dmem_n175), .Y(
        mem_stage_inst_dmem_n133) );
  INV_X1M_A12TS mem_stage_inst_dmem_u34 ( .A(mem_stage_inst_dmem_n175), .Y(
        mem_stage_inst_dmem_n134) );
  INV_X1M_A12TS mem_stage_inst_dmem_u33 ( .A(mem_stage_inst_dmem_n178), .Y(
        mem_stage_inst_dmem_n126) );
  INV_X1M_A12TS mem_stage_inst_dmem_u32 ( .A(mem_stage_inst_dmem_n177), .Y(
        mem_stage_inst_dmem_n127) );
  INV_X1M_A12TS mem_stage_inst_dmem_u31 ( .A(mem_stage_inst_dmem_n177), .Y(
        mem_stage_inst_dmem_n128) );
  INV_X1M_A12TS mem_stage_inst_dmem_u30 ( .A(mem_stage_inst_dmem_n177), .Y(
        mem_stage_inst_dmem_n129) );
  INV_X1M_A12TS mem_stage_inst_dmem_u29 ( .A(mem_stage_inst_dmem_n173), .Y(
        mem_stage_inst_dmem_n140) );
  INV_X1M_A12TS mem_stage_inst_dmem_u28 ( .A(mem_stage_inst_dmem_n173), .Y(
        mem_stage_inst_dmem_n141) );
  INV_X1M_A12TS mem_stage_inst_dmem_u27 ( .A(mem_stage_inst_dmem_n174), .Y(
        mem_stage_inst_dmem_n136) );
  INV_X1M_A12TS mem_stage_inst_dmem_u26 ( .A(mem_stage_inst_dmem_n174), .Y(
        mem_stage_inst_dmem_n137) );
  INV_X1M_A12TS mem_stage_inst_dmem_u25 ( .A(mem_stage_inst_dmem_n174), .Y(
        mem_stage_inst_dmem_n138) );
  INV_X1M_A12TS mem_stage_inst_dmem_u24 ( .A(mem_stage_inst_dmem_n173), .Y(
        mem_stage_inst_dmem_n139) );
  INV_X1M_A12TS mem_stage_inst_dmem_u23 ( .A(mem_stage_inst_dmem_n170), .Y(
        mem_stage_inst_dmem_n150) );
  INV_X1M_A12TS mem_stage_inst_dmem_u22 ( .A(mem_stage_inst_dmem_n169), .Y(
        mem_stage_inst_dmem_n151) );
  INV_X1M_A12TS mem_stage_inst_dmem_u21 ( .A(mem_stage_inst_dmem_n169), .Y(
        mem_stage_inst_dmem_n152) );
  INV_X1M_A12TS mem_stage_inst_dmem_u20 ( .A(mem_stage_inst_dmem_n169), .Y(
        mem_stage_inst_dmem_n153) );
  INV_X1M_A12TS mem_stage_inst_dmem_u19 ( .A(mem_stage_inst_dmem_n168), .Y(
        mem_stage_inst_dmem_n154) );
  INV_X1M_A12TS mem_stage_inst_dmem_u18 ( .A(mem_stage_inst_dmem_n171), .Y(
        mem_stage_inst_dmem_n145) );
  INV_X1M_A12TS mem_stage_inst_dmem_u17 ( .A(mem_stage_inst_dmem_n171), .Y(
        mem_stage_inst_dmem_n146) );
  INV_X1M_A12TS mem_stage_inst_dmem_u16 ( .A(mem_stage_inst_dmem_n171), .Y(
        mem_stage_inst_dmem_n147) );
  INV_X1M_A12TS mem_stage_inst_dmem_u15 ( .A(mem_stage_inst_dmem_n170), .Y(
        mem_stage_inst_dmem_n148) );
  INV_X1M_A12TS mem_stage_inst_dmem_u14 ( .A(mem_stage_inst_dmem_n170), .Y(
        mem_stage_inst_dmem_n149) );
  INV_X1M_A12TS mem_stage_inst_dmem_u13 ( .A(mem_stage_inst_dmem_n167), .Y(
        mem_stage_inst_dmem_n159) );
  INV_X1M_A12TS mem_stage_inst_dmem_u12 ( .A(mem_stage_inst_dmem_n166), .Y(
        mem_stage_inst_dmem_n160) );
  INV_X1M_A12TS mem_stage_inst_dmem_u11 ( .A(mem_stage_inst_dmem_n166), .Y(
        mem_stage_inst_dmem_n161) );
  INV_X1M_A12TS mem_stage_inst_dmem_u10 ( .A(mem_stage_inst_dmem_n166), .Y(
        mem_stage_inst_dmem_n162) );
  INV_X1M_A12TS mem_stage_inst_dmem_u9 ( .A(mem_stage_inst_dmem_n165), .Y(
        mem_stage_inst_dmem_n163) );
  INV_X1M_A12TS mem_stage_inst_dmem_u8 ( .A(mem_stage_inst_dmem_n168), .Y(
        mem_stage_inst_dmem_n155) );
  INV_X1M_A12TS mem_stage_inst_dmem_u7 ( .A(mem_stage_inst_dmem_n168), .Y(
        mem_stage_inst_dmem_n156) );
  INV_X1M_A12TS mem_stage_inst_dmem_u6 ( .A(mem_stage_inst_dmem_n167), .Y(
        mem_stage_inst_dmem_n157) );
  INV_X1M_A12TS mem_stage_inst_dmem_u5 ( .A(mem_stage_inst_dmem_n167), .Y(
        mem_stage_inst_dmem_n158) );
  INV_X1M_A12TS mem_stage_inst_dmem_u4 ( .A(mem_stage_inst_dmem_n172), .Y(
        mem_stage_inst_dmem_n142) );
  INV_X1M_A12TS mem_stage_inst_dmem_u3 ( .A(mem_stage_inst_dmem_n172), .Y(
        mem_stage_inst_dmem_n143) );
  INV_X1M_A12TS mem_stage_inst_dmem_u2 ( .A(mem_stage_inst_dmem_n172), .Y(
        mem_stage_inst_dmem_n144) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__0_ ( .D(
        mem_stage_inst_dmem_n597), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__1_ ( .D(
        mem_stage_inst_dmem_n598), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__2_ ( .D(
        mem_stage_inst_dmem_n599), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__3_ ( .D(
        mem_stage_inst_dmem_n600), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__4_ ( .D(
        mem_stage_inst_dmem_n601), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__5_ ( .D(
        mem_stage_inst_dmem_n602), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__6_ ( .D(
        mem_stage_inst_dmem_n603), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__7_ ( .D(
        mem_stage_inst_dmem_n604), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__8_ ( .D(
        mem_stage_inst_dmem_n605), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__9_ ( .D(
        mem_stage_inst_dmem_n606), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__10_ ( .D(
        mem_stage_inst_dmem_n607), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__11_ ( .D(
        mem_stage_inst_dmem_n608), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__12_ ( .D(
        mem_stage_inst_dmem_n609), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__13_ ( .D(
        mem_stage_inst_dmem_n610), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__14_ ( .D(
        mem_stage_inst_dmem_n611), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_2__15_ ( .D(
        mem_stage_inst_dmem_n612), .CK(clk), .Q(mem_stage_inst_dmem_ram_2__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__0_ ( .D(
        mem_stage_inst_dmem_n661), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__1_ ( .D(
        mem_stage_inst_dmem_n662), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__2_ ( .D(
        mem_stage_inst_dmem_n663), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__3_ ( .D(
        mem_stage_inst_dmem_n664), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__4_ ( .D(
        mem_stage_inst_dmem_n665), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__5_ ( .D(
        mem_stage_inst_dmem_n666), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__6_ ( .D(
        mem_stage_inst_dmem_n667), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__7_ ( .D(
        mem_stage_inst_dmem_n668), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__8_ ( .D(
        mem_stage_inst_dmem_n669), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__9_ ( .D(
        mem_stage_inst_dmem_n670), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__10_ ( .D(
        mem_stage_inst_dmem_n671), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__11_ ( .D(
        mem_stage_inst_dmem_n672), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__12_ ( .D(
        mem_stage_inst_dmem_n673), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__13_ ( .D(
        mem_stage_inst_dmem_n674), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__14_ ( .D(
        mem_stage_inst_dmem_n675), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_6__15_ ( .D(
        mem_stage_inst_dmem_n676), .CK(clk), .Q(mem_stage_inst_dmem_ram_6__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__0_ ( .D(
        mem_stage_inst_dmem_n725), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__1_ ( .D(
        mem_stage_inst_dmem_n726), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__2_ ( .D(
        mem_stage_inst_dmem_n727), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__3_ ( .D(
        mem_stage_inst_dmem_n728), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__4_ ( .D(
        mem_stage_inst_dmem_n729), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__5_ ( .D(
        mem_stage_inst_dmem_n730), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__6_ ( .D(
        mem_stage_inst_dmem_n731), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__7_ ( .D(
        mem_stage_inst_dmem_n732), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__8_ ( .D(
        mem_stage_inst_dmem_n733), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__9_ ( .D(
        mem_stage_inst_dmem_n734), .CK(clk), .Q(mem_stage_inst_dmem_ram_10__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__10_ ( .D(
        mem_stage_inst_dmem_n735), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_10__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__11_ ( .D(
        mem_stage_inst_dmem_n736), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_10__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__12_ ( .D(
        mem_stage_inst_dmem_n737), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_10__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__13_ ( .D(
        mem_stage_inst_dmem_n738), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_10__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__14_ ( .D(
        mem_stage_inst_dmem_n739), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_10__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_10__15_ ( .D(
        mem_stage_inst_dmem_n740), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_10__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__0_ ( .D(
        mem_stage_inst_dmem_n789), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__1_ ( .D(
        mem_stage_inst_dmem_n790), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__2_ ( .D(
        mem_stage_inst_dmem_n791), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__3_ ( .D(
        mem_stage_inst_dmem_n792), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__4_ ( .D(
        mem_stage_inst_dmem_n793), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__5_ ( .D(
        mem_stage_inst_dmem_n794), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__6_ ( .D(
        mem_stage_inst_dmem_n795), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__7_ ( .D(
        mem_stage_inst_dmem_n796), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__8_ ( .D(
        mem_stage_inst_dmem_n797), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__9_ ( .D(
        mem_stage_inst_dmem_n798), .CK(clk), .Q(mem_stage_inst_dmem_ram_14__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__10_ ( .D(
        mem_stage_inst_dmem_n799), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_14__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__11_ ( .D(
        mem_stage_inst_dmem_n800), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_14__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__12_ ( .D(
        mem_stage_inst_dmem_n801), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_14__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__13_ ( .D(
        mem_stage_inst_dmem_n802), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_14__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__14_ ( .D(
        mem_stage_inst_dmem_n803), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_14__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_14__15_ ( .D(
        mem_stage_inst_dmem_n804), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_14__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__0_ ( .D(
        mem_stage_inst_dmem_n853), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__1_ ( .D(
        mem_stage_inst_dmem_n854), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__2_ ( .D(
        mem_stage_inst_dmem_n855), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__3_ ( .D(
        mem_stage_inst_dmem_n856), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__4_ ( .D(
        mem_stage_inst_dmem_n857), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__5_ ( .D(
        mem_stage_inst_dmem_n858), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__6_ ( .D(
        mem_stage_inst_dmem_n859), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__7_ ( .D(
        mem_stage_inst_dmem_n860), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__8_ ( .D(
        mem_stage_inst_dmem_n861), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__9_ ( .D(
        mem_stage_inst_dmem_n862), .CK(clk), .Q(mem_stage_inst_dmem_ram_18__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__10_ ( .D(
        mem_stage_inst_dmem_n863), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_18__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__11_ ( .D(
        mem_stage_inst_dmem_n864), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_18__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__12_ ( .D(
        mem_stage_inst_dmem_n865), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_18__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__13_ ( .D(
        mem_stage_inst_dmem_n866), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_18__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__14_ ( .D(
        mem_stage_inst_dmem_n867), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_18__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_18__15_ ( .D(
        mem_stage_inst_dmem_n868), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_18__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__0_ ( .D(
        mem_stage_inst_dmem_n917), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__1_ ( .D(
        mem_stage_inst_dmem_n918), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__2_ ( .D(
        mem_stage_inst_dmem_n919), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__3_ ( .D(
        mem_stage_inst_dmem_n920), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__4_ ( .D(
        mem_stage_inst_dmem_n921), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__5_ ( .D(
        mem_stage_inst_dmem_n922), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__6_ ( .D(
        mem_stage_inst_dmem_n923), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__7_ ( .D(
        mem_stage_inst_dmem_n924), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__8_ ( .D(
        mem_stage_inst_dmem_n925), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__9_ ( .D(
        mem_stage_inst_dmem_n926), .CK(clk), .Q(mem_stage_inst_dmem_ram_22__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__10_ ( .D(
        mem_stage_inst_dmem_n927), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_22__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__11_ ( .D(
        mem_stage_inst_dmem_n928), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_22__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__12_ ( .D(
        mem_stage_inst_dmem_n929), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_22__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__13_ ( .D(
        mem_stage_inst_dmem_n930), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_22__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__14_ ( .D(
        mem_stage_inst_dmem_n931), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_22__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_22__15_ ( .D(
        mem_stage_inst_dmem_n932), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_22__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__0_ ( .D(
        mem_stage_inst_dmem_n981), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__1_ ( .D(
        mem_stage_inst_dmem_n982), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__2_ ( .D(
        mem_stage_inst_dmem_n983), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__3_ ( .D(
        mem_stage_inst_dmem_n984), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__4_ ( .D(
        mem_stage_inst_dmem_n985), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__5_ ( .D(
        mem_stage_inst_dmem_n986), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__6_ ( .D(
        mem_stage_inst_dmem_n987), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__7_ ( .D(
        mem_stage_inst_dmem_n988), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__8_ ( .D(
        mem_stage_inst_dmem_n989), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__9_ ( .D(
        mem_stage_inst_dmem_n990), .CK(clk), .Q(mem_stage_inst_dmem_ram_26__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__10_ ( .D(
        mem_stage_inst_dmem_n991), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_26__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__11_ ( .D(
        mem_stage_inst_dmem_n992), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_26__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__12_ ( .D(
        mem_stage_inst_dmem_n993), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_26__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__13_ ( .D(
        mem_stage_inst_dmem_n994), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_26__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__14_ ( .D(
        mem_stage_inst_dmem_n995), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_26__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_26__15_ ( .D(
        mem_stage_inst_dmem_n996), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_26__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__0_ ( .D(
        mem_stage_inst_dmem_n1045), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__1_ ( .D(
        mem_stage_inst_dmem_n1046), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__2_ ( .D(
        mem_stage_inst_dmem_n1047), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__3_ ( .D(
        mem_stage_inst_dmem_n1048), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__4_ ( .D(
        mem_stage_inst_dmem_n1049), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__5_ ( .D(
        mem_stage_inst_dmem_n1050), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__6_ ( .D(
        mem_stage_inst_dmem_n1051), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__7_ ( .D(
        mem_stage_inst_dmem_n1052), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__8_ ( .D(
        mem_stage_inst_dmem_n1053), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__9_ ( .D(
        mem_stage_inst_dmem_n1054), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__10_ ( .D(
        mem_stage_inst_dmem_n1055), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__11_ ( .D(
        mem_stage_inst_dmem_n1056), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__12_ ( .D(
        mem_stage_inst_dmem_n1057), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__13_ ( .D(
        mem_stage_inst_dmem_n1058), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__14_ ( .D(
        mem_stage_inst_dmem_n1059), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_30__15_ ( .D(
        mem_stage_inst_dmem_n1060), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_30__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__0_ ( .D(
        mem_stage_inst_dmem_n1109), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__1_ ( .D(
        mem_stage_inst_dmem_n1110), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__2_ ( .D(
        mem_stage_inst_dmem_n1111), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__3_ ( .D(
        mem_stage_inst_dmem_n1112), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__4_ ( .D(
        mem_stage_inst_dmem_n1113), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__5_ ( .D(
        mem_stage_inst_dmem_n1114), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__6_ ( .D(
        mem_stage_inst_dmem_n1115), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__7_ ( .D(
        mem_stage_inst_dmem_n1116), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__8_ ( .D(
        mem_stage_inst_dmem_n1117), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__9_ ( .D(
        mem_stage_inst_dmem_n1118), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__10_ ( .D(
        mem_stage_inst_dmem_n1119), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__11_ ( .D(
        mem_stage_inst_dmem_n1120), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__12_ ( .D(
        mem_stage_inst_dmem_n1121), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__13_ ( .D(
        mem_stage_inst_dmem_n1122), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__14_ ( .D(
        mem_stage_inst_dmem_n1123), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_34__15_ ( .D(
        mem_stage_inst_dmem_n1124), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_34__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__0_ ( .D(
        mem_stage_inst_dmem_n1173), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__1_ ( .D(
        mem_stage_inst_dmem_n1174), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__2_ ( .D(
        mem_stage_inst_dmem_n1175), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__3_ ( .D(
        mem_stage_inst_dmem_n1176), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__4_ ( .D(
        mem_stage_inst_dmem_n1177), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__5_ ( .D(
        mem_stage_inst_dmem_n1178), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__6_ ( .D(
        mem_stage_inst_dmem_n1179), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__7_ ( .D(
        mem_stage_inst_dmem_n1180), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__8_ ( .D(
        mem_stage_inst_dmem_n1181), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__9_ ( .D(
        mem_stage_inst_dmem_n1182), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__10_ ( .D(
        mem_stage_inst_dmem_n1183), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__11_ ( .D(
        mem_stage_inst_dmem_n1184), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__12_ ( .D(
        mem_stage_inst_dmem_n1185), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__13_ ( .D(
        mem_stage_inst_dmem_n1186), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__14_ ( .D(
        mem_stage_inst_dmem_n1187), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_38__15_ ( .D(
        mem_stage_inst_dmem_n1188), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_38__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__0_ ( .D(
        mem_stage_inst_dmem_n1237), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__1_ ( .D(
        mem_stage_inst_dmem_n1238), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__2_ ( .D(
        mem_stage_inst_dmem_n1239), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__3_ ( .D(
        mem_stage_inst_dmem_n1240), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__4_ ( .D(
        mem_stage_inst_dmem_n1241), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__5_ ( .D(
        mem_stage_inst_dmem_n1242), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__6_ ( .D(
        mem_stage_inst_dmem_n1243), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__7_ ( .D(
        mem_stage_inst_dmem_n1244), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__8_ ( .D(
        mem_stage_inst_dmem_n1245), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__9_ ( .D(
        mem_stage_inst_dmem_n1246), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__10_ ( .D(
        mem_stage_inst_dmem_n1247), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__11_ ( .D(
        mem_stage_inst_dmem_n1248), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__12_ ( .D(
        mem_stage_inst_dmem_n1249), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__13_ ( .D(
        mem_stage_inst_dmem_n1250), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__14_ ( .D(
        mem_stage_inst_dmem_n1251), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_42__15_ ( .D(
        mem_stage_inst_dmem_n1252), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_42__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__0_ ( .D(
        mem_stage_inst_dmem_n1301), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__1_ ( .D(
        mem_stage_inst_dmem_n1302), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__2_ ( .D(
        mem_stage_inst_dmem_n1303), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__3_ ( .D(
        mem_stage_inst_dmem_n1304), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__4_ ( .D(
        mem_stage_inst_dmem_n1305), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__5_ ( .D(
        mem_stage_inst_dmem_n1306), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__6_ ( .D(
        mem_stage_inst_dmem_n1307), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__7_ ( .D(
        mem_stage_inst_dmem_n1308), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__8_ ( .D(
        mem_stage_inst_dmem_n1309), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__9_ ( .D(
        mem_stage_inst_dmem_n1310), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__10_ ( .D(
        mem_stage_inst_dmem_n1311), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__11_ ( .D(
        mem_stage_inst_dmem_n1312), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__12_ ( .D(
        mem_stage_inst_dmem_n1313), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__13_ ( .D(
        mem_stage_inst_dmem_n1314), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__14_ ( .D(
        mem_stage_inst_dmem_n1315), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_46__15_ ( .D(
        mem_stage_inst_dmem_n1316), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_46__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__0_ ( .D(
        mem_stage_inst_dmem_n1365), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__1_ ( .D(
        mem_stage_inst_dmem_n1366), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__2_ ( .D(
        mem_stage_inst_dmem_n1367), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__3_ ( .D(
        mem_stage_inst_dmem_n1368), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__4_ ( .D(
        mem_stage_inst_dmem_n1369), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__5_ ( .D(
        mem_stage_inst_dmem_n1370), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__6_ ( .D(
        mem_stage_inst_dmem_n1371), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__7_ ( .D(
        mem_stage_inst_dmem_n1372), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__8_ ( .D(
        mem_stage_inst_dmem_n1373), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__9_ ( .D(
        mem_stage_inst_dmem_n1374), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__10_ ( .D(
        mem_stage_inst_dmem_n1375), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__11_ ( .D(
        mem_stage_inst_dmem_n1376), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__12_ ( .D(
        mem_stage_inst_dmem_n1377), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__13_ ( .D(
        mem_stage_inst_dmem_n1378), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__14_ ( .D(
        mem_stage_inst_dmem_n1379), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_50__15_ ( .D(
        mem_stage_inst_dmem_n1380), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_50__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__0_ ( .D(
        mem_stage_inst_dmem_n1429), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__1_ ( .D(
        mem_stage_inst_dmem_n1430), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__2_ ( .D(
        mem_stage_inst_dmem_n1431), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__3_ ( .D(
        mem_stage_inst_dmem_n1432), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__4_ ( .D(
        mem_stage_inst_dmem_n1433), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__5_ ( .D(
        mem_stage_inst_dmem_n1434), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__6_ ( .D(
        mem_stage_inst_dmem_n1435), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__7_ ( .D(
        mem_stage_inst_dmem_n1436), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__8_ ( .D(
        mem_stage_inst_dmem_n1437), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__9_ ( .D(
        mem_stage_inst_dmem_n1438), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__10_ ( .D(
        mem_stage_inst_dmem_n1439), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__11_ ( .D(
        mem_stage_inst_dmem_n1440), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__12_ ( .D(
        mem_stage_inst_dmem_n1441), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__13_ ( .D(
        mem_stage_inst_dmem_n1442), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__14_ ( .D(
        mem_stage_inst_dmem_n1443), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_54__15_ ( .D(
        mem_stage_inst_dmem_n1444), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_54__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__0_ ( .D(
        mem_stage_inst_dmem_n1493), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__1_ ( .D(
        mem_stage_inst_dmem_n1494), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__2_ ( .D(
        mem_stage_inst_dmem_n1495), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__3_ ( .D(
        mem_stage_inst_dmem_n1496), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__4_ ( .D(
        mem_stage_inst_dmem_n1497), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__5_ ( .D(
        mem_stage_inst_dmem_n1498), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__6_ ( .D(
        mem_stage_inst_dmem_n1499), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__7_ ( .D(
        mem_stage_inst_dmem_n1500), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__8_ ( .D(
        mem_stage_inst_dmem_n1501), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__9_ ( .D(
        mem_stage_inst_dmem_n1502), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__10_ ( .D(
        mem_stage_inst_dmem_n1503), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__11_ ( .D(
        mem_stage_inst_dmem_n1504), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__12_ ( .D(
        mem_stage_inst_dmem_n1505), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__13_ ( .D(
        mem_stage_inst_dmem_n1506), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__14_ ( .D(
        mem_stage_inst_dmem_n1507), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_58__15_ ( .D(
        mem_stage_inst_dmem_n1508), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_58__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__0_ ( .D(
        mem_stage_inst_dmem_n1557), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__1_ ( .D(
        mem_stage_inst_dmem_n1558), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__2_ ( .D(
        mem_stage_inst_dmem_n1559), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__3_ ( .D(
        mem_stage_inst_dmem_n1560), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__4_ ( .D(
        mem_stage_inst_dmem_n1561), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__5_ ( .D(
        mem_stage_inst_dmem_n1562), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__6_ ( .D(
        mem_stage_inst_dmem_n1563), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__7_ ( .D(
        mem_stage_inst_dmem_n1564), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__8_ ( .D(
        mem_stage_inst_dmem_n1565), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__9_ ( .D(
        mem_stage_inst_dmem_n1566), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__10_ ( .D(
        mem_stage_inst_dmem_n1567), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__11_ ( .D(
        mem_stage_inst_dmem_n1568), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__12_ ( .D(
        mem_stage_inst_dmem_n1569), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__13_ ( .D(
        mem_stage_inst_dmem_n1570), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__14_ ( .D(
        mem_stage_inst_dmem_n1571), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_62__15_ ( .D(
        mem_stage_inst_dmem_n1572), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_62__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__0_ ( .D(
        mem_stage_inst_dmem_n1621), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__1_ ( .D(
        mem_stage_inst_dmem_n1622), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__2_ ( .D(
        mem_stage_inst_dmem_n1623), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__3_ ( .D(
        mem_stage_inst_dmem_n1624), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__4_ ( .D(
        mem_stage_inst_dmem_n1625), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__5_ ( .D(
        mem_stage_inst_dmem_n1626), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__6_ ( .D(
        mem_stage_inst_dmem_n1627), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__7_ ( .D(
        mem_stage_inst_dmem_n1628), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__8_ ( .D(
        mem_stage_inst_dmem_n1629), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__9_ ( .D(
        mem_stage_inst_dmem_n1630), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__10_ ( .D(
        mem_stage_inst_dmem_n1631), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__11_ ( .D(
        mem_stage_inst_dmem_n1632), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__12_ ( .D(
        mem_stage_inst_dmem_n1633), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__13_ ( .D(
        mem_stage_inst_dmem_n1634), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__14_ ( .D(
        mem_stage_inst_dmem_n1635), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_66__15_ ( .D(
        mem_stage_inst_dmem_n1636), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_66__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__0_ ( .D(
        mem_stage_inst_dmem_n1685), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__1_ ( .D(
        mem_stage_inst_dmem_n1686), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__2_ ( .D(
        mem_stage_inst_dmem_n1687), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__3_ ( .D(
        mem_stage_inst_dmem_n1688), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__4_ ( .D(
        mem_stage_inst_dmem_n1689), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__5_ ( .D(
        mem_stage_inst_dmem_n1690), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__6_ ( .D(
        mem_stage_inst_dmem_n1691), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__7_ ( .D(
        mem_stage_inst_dmem_n1692), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__8_ ( .D(
        mem_stage_inst_dmem_n1693), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__9_ ( .D(
        mem_stage_inst_dmem_n1694), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__10_ ( .D(
        mem_stage_inst_dmem_n1695), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__11_ ( .D(
        mem_stage_inst_dmem_n1696), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__12_ ( .D(
        mem_stage_inst_dmem_n1697), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__13_ ( .D(
        mem_stage_inst_dmem_n1698), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__14_ ( .D(
        mem_stage_inst_dmem_n1699), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_70__15_ ( .D(
        mem_stage_inst_dmem_n1700), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_70__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__0_ ( .D(
        mem_stage_inst_dmem_n1749), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__1_ ( .D(
        mem_stage_inst_dmem_n1750), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__2_ ( .D(
        mem_stage_inst_dmem_n1751), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__3_ ( .D(
        mem_stage_inst_dmem_n1752), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__4_ ( .D(
        mem_stage_inst_dmem_n1753), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__5_ ( .D(
        mem_stage_inst_dmem_n1754), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__6_ ( .D(
        mem_stage_inst_dmem_n1755), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__7_ ( .D(
        mem_stage_inst_dmem_n1756), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__8_ ( .D(
        mem_stage_inst_dmem_n1757), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__9_ ( .D(
        mem_stage_inst_dmem_n1758), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__10_ ( .D(
        mem_stage_inst_dmem_n1759), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__11_ ( .D(
        mem_stage_inst_dmem_n1760), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__12_ ( .D(
        mem_stage_inst_dmem_n1761), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__13_ ( .D(
        mem_stage_inst_dmem_n1762), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__14_ ( .D(
        mem_stage_inst_dmem_n1763), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_74__15_ ( .D(
        mem_stage_inst_dmem_n1764), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_74__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__0_ ( .D(
        mem_stage_inst_dmem_n1813), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__1_ ( .D(
        mem_stage_inst_dmem_n1814), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__2_ ( .D(
        mem_stage_inst_dmem_n1815), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__3_ ( .D(
        mem_stage_inst_dmem_n1816), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__4_ ( .D(
        mem_stage_inst_dmem_n1817), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__5_ ( .D(
        mem_stage_inst_dmem_n1818), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__6_ ( .D(
        mem_stage_inst_dmem_n1819), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__7_ ( .D(
        mem_stage_inst_dmem_n1820), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__8_ ( .D(
        mem_stage_inst_dmem_n1821), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__9_ ( .D(
        mem_stage_inst_dmem_n1822), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__10_ ( .D(
        mem_stage_inst_dmem_n1823), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__11_ ( .D(
        mem_stage_inst_dmem_n1824), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__12_ ( .D(
        mem_stage_inst_dmem_n1825), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__13_ ( .D(
        mem_stage_inst_dmem_n1826), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__14_ ( .D(
        mem_stage_inst_dmem_n1827), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_78__15_ ( .D(
        mem_stage_inst_dmem_n1828), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_78__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__0_ ( .D(
        mem_stage_inst_dmem_n1877), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__1_ ( .D(
        mem_stage_inst_dmem_n1878), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__2_ ( .D(
        mem_stage_inst_dmem_n1879), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__3_ ( .D(
        mem_stage_inst_dmem_n1880), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__4_ ( .D(
        mem_stage_inst_dmem_n1881), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__5_ ( .D(
        mem_stage_inst_dmem_n1882), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__6_ ( .D(
        mem_stage_inst_dmem_n1883), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__7_ ( .D(
        mem_stage_inst_dmem_n1884), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__8_ ( .D(
        mem_stage_inst_dmem_n1885), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__9_ ( .D(
        mem_stage_inst_dmem_n1886), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__10_ ( .D(
        mem_stage_inst_dmem_n1887), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__11_ ( .D(
        mem_stage_inst_dmem_n1888), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__12_ ( .D(
        mem_stage_inst_dmem_n1889), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__13_ ( .D(
        mem_stage_inst_dmem_n1890), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__14_ ( .D(
        mem_stage_inst_dmem_n1891), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_82__15_ ( .D(
        mem_stage_inst_dmem_n1892), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_82__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__0_ ( .D(
        mem_stage_inst_dmem_n1941), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__1_ ( .D(
        mem_stage_inst_dmem_n1942), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__2_ ( .D(
        mem_stage_inst_dmem_n1943), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__3_ ( .D(
        mem_stage_inst_dmem_n1944), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__4_ ( .D(
        mem_stage_inst_dmem_n1945), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__5_ ( .D(
        mem_stage_inst_dmem_n1946), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__6_ ( .D(
        mem_stage_inst_dmem_n1947), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__7_ ( .D(
        mem_stage_inst_dmem_n1948), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__8_ ( .D(
        mem_stage_inst_dmem_n1949), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__9_ ( .D(
        mem_stage_inst_dmem_n1950), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__10_ ( .D(
        mem_stage_inst_dmem_n1951), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__11_ ( .D(
        mem_stage_inst_dmem_n1952), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__12_ ( .D(
        mem_stage_inst_dmem_n1953), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__13_ ( .D(
        mem_stage_inst_dmem_n1954), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__14_ ( .D(
        mem_stage_inst_dmem_n1955), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_86__15_ ( .D(
        mem_stage_inst_dmem_n1956), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_86__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__0_ ( .D(
        mem_stage_inst_dmem_n2005), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__1_ ( .D(
        mem_stage_inst_dmem_n2006), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__2_ ( .D(
        mem_stage_inst_dmem_n2007), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__3_ ( .D(
        mem_stage_inst_dmem_n2008), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__4_ ( .D(
        mem_stage_inst_dmem_n2009), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__5_ ( .D(
        mem_stage_inst_dmem_n2010), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__6_ ( .D(
        mem_stage_inst_dmem_n2011), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__7_ ( .D(
        mem_stage_inst_dmem_n2012), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__8_ ( .D(
        mem_stage_inst_dmem_n2013), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__9_ ( .D(
        mem_stage_inst_dmem_n2014), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__10_ ( .D(
        mem_stage_inst_dmem_n2015), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__11_ ( .D(
        mem_stage_inst_dmem_n2016), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__12_ ( .D(
        mem_stage_inst_dmem_n2017), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__13_ ( .D(
        mem_stage_inst_dmem_n2018), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__14_ ( .D(
        mem_stage_inst_dmem_n2019), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_90__15_ ( .D(
        mem_stage_inst_dmem_n2020), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_90__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__0_ ( .D(
        mem_stage_inst_dmem_n2069), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__1_ ( .D(
        mem_stage_inst_dmem_n2070), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__2_ ( .D(
        mem_stage_inst_dmem_n2071), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__3_ ( .D(
        mem_stage_inst_dmem_n2072), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__4_ ( .D(
        mem_stage_inst_dmem_n2073), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__5_ ( .D(
        mem_stage_inst_dmem_n2074), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__6_ ( .D(
        mem_stage_inst_dmem_n2075), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__7_ ( .D(
        mem_stage_inst_dmem_n2076), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__8_ ( .D(
        mem_stage_inst_dmem_n2077), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__9_ ( .D(
        mem_stage_inst_dmem_n2078), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__10_ ( .D(
        mem_stage_inst_dmem_n2079), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__11_ ( .D(
        mem_stage_inst_dmem_n2080), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__12_ ( .D(
        mem_stage_inst_dmem_n2081), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__13_ ( .D(
        mem_stage_inst_dmem_n2082), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__14_ ( .D(
        mem_stage_inst_dmem_n2083), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_94__15_ ( .D(
        mem_stage_inst_dmem_n2084), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_94__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__0_ ( .D(
        mem_stage_inst_dmem_n2133), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__1_ ( .D(
        mem_stage_inst_dmem_n2134), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__2_ ( .D(
        mem_stage_inst_dmem_n2135), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__3_ ( .D(
        mem_stage_inst_dmem_n2136), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__4_ ( .D(
        mem_stage_inst_dmem_n2137), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__5_ ( .D(
        mem_stage_inst_dmem_n2138), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__6_ ( .D(
        mem_stage_inst_dmem_n2139), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__7_ ( .D(
        mem_stage_inst_dmem_n2140), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__8_ ( .D(
        mem_stage_inst_dmem_n2141), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__9_ ( .D(
        mem_stage_inst_dmem_n2142), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__10_ ( .D(
        mem_stage_inst_dmem_n2143), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__11_ ( .D(
        mem_stage_inst_dmem_n2144), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__12_ ( .D(
        mem_stage_inst_dmem_n2145), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__13_ ( .D(
        mem_stage_inst_dmem_n2146), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__14_ ( .D(
        mem_stage_inst_dmem_n2147), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_98__15_ ( .D(
        mem_stage_inst_dmem_n2148), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_98__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__0_ ( .D(
        mem_stage_inst_dmem_n2197), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__1_ ( .D(
        mem_stage_inst_dmem_n2198), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__2_ ( .D(
        mem_stage_inst_dmem_n2199), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__3_ ( .D(
        mem_stage_inst_dmem_n2200), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__4_ ( .D(
        mem_stage_inst_dmem_n2201), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__5_ ( .D(
        mem_stage_inst_dmem_n2202), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__6_ ( .D(
        mem_stage_inst_dmem_n2203), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__7_ ( .D(
        mem_stage_inst_dmem_n2204), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__8_ ( .D(
        mem_stage_inst_dmem_n2205), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__9_ ( .D(
        mem_stage_inst_dmem_n2206), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__10_ ( .D(
        mem_stage_inst_dmem_n2207), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__11_ ( .D(
        mem_stage_inst_dmem_n2208), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__12_ ( .D(
        mem_stage_inst_dmem_n2209), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__13_ ( .D(
        mem_stage_inst_dmem_n2210), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__14_ ( .D(
        mem_stage_inst_dmem_n2211), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_102__15_ ( .D(
        mem_stage_inst_dmem_n2212), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_102__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__0_ ( .D(
        mem_stage_inst_dmem_n2261), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__1_ ( .D(
        mem_stage_inst_dmem_n2262), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__2_ ( .D(
        mem_stage_inst_dmem_n2263), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__3_ ( .D(
        mem_stage_inst_dmem_n2264), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__4_ ( .D(
        mem_stage_inst_dmem_n2265), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__5_ ( .D(
        mem_stage_inst_dmem_n2266), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__6_ ( .D(
        mem_stage_inst_dmem_n2267), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__7_ ( .D(
        mem_stage_inst_dmem_n2268), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__8_ ( .D(
        mem_stage_inst_dmem_n2269), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__9_ ( .D(
        mem_stage_inst_dmem_n2270), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__10_ ( .D(
        mem_stage_inst_dmem_n2271), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__11_ ( .D(
        mem_stage_inst_dmem_n2272), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__12_ ( .D(
        mem_stage_inst_dmem_n2273), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__13_ ( .D(
        mem_stage_inst_dmem_n2274), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__14_ ( .D(
        mem_stage_inst_dmem_n2275), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_106__15_ ( .D(
        mem_stage_inst_dmem_n2276), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_106__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__0_ ( .D(
        mem_stage_inst_dmem_n2325), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__1_ ( .D(
        mem_stage_inst_dmem_n2326), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__2_ ( .D(
        mem_stage_inst_dmem_n2327), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__3_ ( .D(
        mem_stage_inst_dmem_n2328), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__4_ ( .D(
        mem_stage_inst_dmem_n2329), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__5_ ( .D(
        mem_stage_inst_dmem_n2330), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__6_ ( .D(
        mem_stage_inst_dmem_n2331), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__7_ ( .D(
        mem_stage_inst_dmem_n2332), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__8_ ( .D(
        mem_stage_inst_dmem_n2333), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__9_ ( .D(
        mem_stage_inst_dmem_n2334), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__10_ ( .D(
        mem_stage_inst_dmem_n2335), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__11_ ( .D(
        mem_stage_inst_dmem_n2336), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__12_ ( .D(
        mem_stage_inst_dmem_n2337), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__13_ ( .D(
        mem_stage_inst_dmem_n2338), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__14_ ( .D(
        mem_stage_inst_dmem_n2339), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_110__15_ ( .D(
        mem_stage_inst_dmem_n2340), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_110__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__0_ ( .D(
        mem_stage_inst_dmem_n2389), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__1_ ( .D(
        mem_stage_inst_dmem_n2390), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__2_ ( .D(
        mem_stage_inst_dmem_n2391), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__3_ ( .D(
        mem_stage_inst_dmem_n2392), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__4_ ( .D(
        mem_stage_inst_dmem_n2393), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__5_ ( .D(
        mem_stage_inst_dmem_n2394), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__6_ ( .D(
        mem_stage_inst_dmem_n2395), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__7_ ( .D(
        mem_stage_inst_dmem_n2396), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__8_ ( .D(
        mem_stage_inst_dmem_n2397), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__9_ ( .D(
        mem_stage_inst_dmem_n2398), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__10_ ( .D(
        mem_stage_inst_dmem_n2399), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__11_ ( .D(
        mem_stage_inst_dmem_n2400), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__12_ ( .D(
        mem_stage_inst_dmem_n2401), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__13_ ( .D(
        mem_stage_inst_dmem_n2402), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__14_ ( .D(
        mem_stage_inst_dmem_n2403), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_114__15_ ( .D(
        mem_stage_inst_dmem_n2404), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_114__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__0_ ( .D(
        mem_stage_inst_dmem_n2453), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__1_ ( .D(
        mem_stage_inst_dmem_n2454), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__2_ ( .D(
        mem_stage_inst_dmem_n2455), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__3_ ( .D(
        mem_stage_inst_dmem_n2456), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__4_ ( .D(
        mem_stage_inst_dmem_n2457), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__5_ ( .D(
        mem_stage_inst_dmem_n2458), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__6_ ( .D(
        mem_stage_inst_dmem_n2459), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__7_ ( .D(
        mem_stage_inst_dmem_n2460), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__8_ ( .D(
        mem_stage_inst_dmem_n2461), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__9_ ( .D(
        mem_stage_inst_dmem_n2462), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__10_ ( .D(
        mem_stage_inst_dmem_n2463), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__11_ ( .D(
        mem_stage_inst_dmem_n2464), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__12_ ( .D(
        mem_stage_inst_dmem_n2465), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__13_ ( .D(
        mem_stage_inst_dmem_n2466), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__14_ ( .D(
        mem_stage_inst_dmem_n2467), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_118__15_ ( .D(
        mem_stage_inst_dmem_n2468), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_118__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__0_ ( .D(
        mem_stage_inst_dmem_n2517), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__1_ ( .D(
        mem_stage_inst_dmem_n2518), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__2_ ( .D(
        mem_stage_inst_dmem_n2519), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__3_ ( .D(
        mem_stage_inst_dmem_n2520), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__4_ ( .D(
        mem_stage_inst_dmem_n2521), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__5_ ( .D(
        mem_stage_inst_dmem_n2522), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__6_ ( .D(
        mem_stage_inst_dmem_n2523), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__7_ ( .D(
        mem_stage_inst_dmem_n2524), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__8_ ( .D(
        mem_stage_inst_dmem_n2525), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__9_ ( .D(
        mem_stage_inst_dmem_n2526), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__10_ ( .D(
        mem_stage_inst_dmem_n2527), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__11_ ( .D(
        mem_stage_inst_dmem_n2528), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__12_ ( .D(
        mem_stage_inst_dmem_n2529), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__13_ ( .D(
        mem_stage_inst_dmem_n2530), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__14_ ( .D(
        mem_stage_inst_dmem_n2531), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_122__15_ ( .D(
        mem_stage_inst_dmem_n2532), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_122__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__0_ ( .D(
        mem_stage_inst_dmem_n2581), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__1_ ( .D(
        mem_stage_inst_dmem_n2582), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__2_ ( .D(
        mem_stage_inst_dmem_n2583), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__3_ ( .D(
        mem_stage_inst_dmem_n2584), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__4_ ( .D(
        mem_stage_inst_dmem_n2585), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__5_ ( .D(
        mem_stage_inst_dmem_n2586), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__6_ ( .D(
        mem_stage_inst_dmem_n2587), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__7_ ( .D(
        mem_stage_inst_dmem_n2588), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__8_ ( .D(
        mem_stage_inst_dmem_n2589), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__9_ ( .D(
        mem_stage_inst_dmem_n2590), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__10_ ( .D(
        mem_stage_inst_dmem_n2591), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__11_ ( .D(
        mem_stage_inst_dmem_n2592), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__12_ ( .D(
        mem_stage_inst_dmem_n2593), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__13_ ( .D(
        mem_stage_inst_dmem_n2594), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__14_ ( .D(
        mem_stage_inst_dmem_n2595), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_126__15_ ( .D(
        mem_stage_inst_dmem_n2596), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_126__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__0_ ( .D(
        mem_stage_inst_dmem_n2645), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__1_ ( .D(
        mem_stage_inst_dmem_n2646), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__2_ ( .D(
        mem_stage_inst_dmem_n2647), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__3_ ( .D(
        mem_stage_inst_dmem_n2648), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__4_ ( .D(
        mem_stage_inst_dmem_n2649), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__5_ ( .D(
        mem_stage_inst_dmem_n2650), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__6_ ( .D(
        mem_stage_inst_dmem_n2651), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__7_ ( .D(
        mem_stage_inst_dmem_n2652), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__8_ ( .D(
        mem_stage_inst_dmem_n2653), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__9_ ( .D(
        mem_stage_inst_dmem_n2654), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__10_ ( .D(
        mem_stage_inst_dmem_n2655), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__11_ ( .D(
        mem_stage_inst_dmem_n2656), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__12_ ( .D(
        mem_stage_inst_dmem_n2657), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__13_ ( .D(
        mem_stage_inst_dmem_n2658), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__14_ ( .D(
        mem_stage_inst_dmem_n2659), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_130__15_ ( .D(
        mem_stage_inst_dmem_n2660), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_130__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__0_ ( .D(
        mem_stage_inst_dmem_n2709), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__1_ ( .D(
        mem_stage_inst_dmem_n2710), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__2_ ( .D(
        mem_stage_inst_dmem_n2711), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__3_ ( .D(
        mem_stage_inst_dmem_n2712), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__4_ ( .D(
        mem_stage_inst_dmem_n2713), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__5_ ( .D(
        mem_stage_inst_dmem_n2714), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__6_ ( .D(
        mem_stage_inst_dmem_n2715), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__7_ ( .D(
        mem_stage_inst_dmem_n2716), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__8_ ( .D(
        mem_stage_inst_dmem_n2717), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__9_ ( .D(
        mem_stage_inst_dmem_n2718), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__10_ ( .D(
        mem_stage_inst_dmem_n2719), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__11_ ( .D(
        mem_stage_inst_dmem_n2720), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__12_ ( .D(
        mem_stage_inst_dmem_n2721), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__13_ ( .D(
        mem_stage_inst_dmem_n2722), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__14_ ( .D(
        mem_stage_inst_dmem_n2723), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_134__15_ ( .D(
        mem_stage_inst_dmem_n2724), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_134__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__0_ ( .D(
        mem_stage_inst_dmem_n2773), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__1_ ( .D(
        mem_stage_inst_dmem_n2774), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__2_ ( .D(
        mem_stage_inst_dmem_n2775), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__3_ ( .D(
        mem_stage_inst_dmem_n2776), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__4_ ( .D(
        mem_stage_inst_dmem_n2777), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__5_ ( .D(
        mem_stage_inst_dmem_n2778), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__6_ ( .D(
        mem_stage_inst_dmem_n2779), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__7_ ( .D(
        mem_stage_inst_dmem_n2780), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__8_ ( .D(
        mem_stage_inst_dmem_n2781), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__9_ ( .D(
        mem_stage_inst_dmem_n2782), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__10_ ( .D(
        mem_stage_inst_dmem_n2783), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__11_ ( .D(
        mem_stage_inst_dmem_n2784), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__12_ ( .D(
        mem_stage_inst_dmem_n2785), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__13_ ( .D(
        mem_stage_inst_dmem_n2786), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__14_ ( .D(
        mem_stage_inst_dmem_n2787), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_138__15_ ( .D(
        mem_stage_inst_dmem_n2788), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_138__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__0_ ( .D(
        mem_stage_inst_dmem_n2837), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__1_ ( .D(
        mem_stage_inst_dmem_n2838), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__2_ ( .D(
        mem_stage_inst_dmem_n2839), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__3_ ( .D(
        mem_stage_inst_dmem_n2840), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__4_ ( .D(
        mem_stage_inst_dmem_n2841), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__5_ ( .D(
        mem_stage_inst_dmem_n2842), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__6_ ( .D(
        mem_stage_inst_dmem_n2843), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__7_ ( .D(
        mem_stage_inst_dmem_n2844), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__8_ ( .D(
        mem_stage_inst_dmem_n2845), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__9_ ( .D(
        mem_stage_inst_dmem_n2846), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__10_ ( .D(
        mem_stage_inst_dmem_n2847), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__11_ ( .D(
        mem_stage_inst_dmem_n2848), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__12_ ( .D(
        mem_stage_inst_dmem_n2849), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__13_ ( .D(
        mem_stage_inst_dmem_n2850), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__14_ ( .D(
        mem_stage_inst_dmem_n2851), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_142__15_ ( .D(
        mem_stage_inst_dmem_n2852), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_142__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__0_ ( .D(
        mem_stage_inst_dmem_n2901), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__1_ ( .D(
        mem_stage_inst_dmem_n2902), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__2_ ( .D(
        mem_stage_inst_dmem_n2903), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__3_ ( .D(
        mem_stage_inst_dmem_n2904), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__4_ ( .D(
        mem_stage_inst_dmem_n2905), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__5_ ( .D(
        mem_stage_inst_dmem_n2906), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__6_ ( .D(
        mem_stage_inst_dmem_n2907), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__7_ ( .D(
        mem_stage_inst_dmem_n2908), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__8_ ( .D(
        mem_stage_inst_dmem_n2909), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__9_ ( .D(
        mem_stage_inst_dmem_n2910), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__10_ ( .D(
        mem_stage_inst_dmem_n2911), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__11_ ( .D(
        mem_stage_inst_dmem_n2912), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__12_ ( .D(
        mem_stage_inst_dmem_n2913), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__13_ ( .D(
        mem_stage_inst_dmem_n2914), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__14_ ( .D(
        mem_stage_inst_dmem_n2915), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_146__15_ ( .D(
        mem_stage_inst_dmem_n2916), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_146__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__0_ ( .D(
        mem_stage_inst_dmem_n2965), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__1_ ( .D(
        mem_stage_inst_dmem_n2966), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__2_ ( .D(
        mem_stage_inst_dmem_n2967), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__3_ ( .D(
        mem_stage_inst_dmem_n2968), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__4_ ( .D(
        mem_stage_inst_dmem_n2969), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__5_ ( .D(
        mem_stage_inst_dmem_n2970), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__6_ ( .D(
        mem_stage_inst_dmem_n2971), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__7_ ( .D(
        mem_stage_inst_dmem_n2972), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__8_ ( .D(
        mem_stage_inst_dmem_n2973), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__9_ ( .D(
        mem_stage_inst_dmem_n2974), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__10_ ( .D(
        mem_stage_inst_dmem_n2975), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__11_ ( .D(
        mem_stage_inst_dmem_n2976), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__12_ ( .D(
        mem_stage_inst_dmem_n2977), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__13_ ( .D(
        mem_stage_inst_dmem_n2978), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__14_ ( .D(
        mem_stage_inst_dmem_n2979), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_150__15_ ( .D(
        mem_stage_inst_dmem_n2980), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_150__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__0_ ( .D(
        mem_stage_inst_dmem_n3029), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__1_ ( .D(
        mem_stage_inst_dmem_n3030), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__2_ ( .D(
        mem_stage_inst_dmem_n3031), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__3_ ( .D(
        mem_stage_inst_dmem_n3032), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__4_ ( .D(
        mem_stage_inst_dmem_n3033), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__5_ ( .D(
        mem_stage_inst_dmem_n3034), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__6_ ( .D(
        mem_stage_inst_dmem_n3035), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__7_ ( .D(
        mem_stage_inst_dmem_n3036), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__8_ ( .D(
        mem_stage_inst_dmem_n3037), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__9_ ( .D(
        mem_stage_inst_dmem_n3038), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__10_ ( .D(
        mem_stage_inst_dmem_n3039), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__11_ ( .D(
        mem_stage_inst_dmem_n3040), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__12_ ( .D(
        mem_stage_inst_dmem_n3041), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__13_ ( .D(
        mem_stage_inst_dmem_n3042), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__14_ ( .D(
        mem_stage_inst_dmem_n3043), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_154__15_ ( .D(
        mem_stage_inst_dmem_n3044), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_154__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__0_ ( .D(
        mem_stage_inst_dmem_n3093), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__1_ ( .D(
        mem_stage_inst_dmem_n3094), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__2_ ( .D(
        mem_stage_inst_dmem_n3095), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__3_ ( .D(
        mem_stage_inst_dmem_n3096), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__4_ ( .D(
        mem_stage_inst_dmem_n3097), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__5_ ( .D(
        mem_stage_inst_dmem_n3098), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__6_ ( .D(
        mem_stage_inst_dmem_n3099), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__7_ ( .D(
        mem_stage_inst_dmem_n3100), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__8_ ( .D(
        mem_stage_inst_dmem_n3101), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__9_ ( .D(
        mem_stage_inst_dmem_n3102), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__10_ ( .D(
        mem_stage_inst_dmem_n3103), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__11_ ( .D(
        mem_stage_inst_dmem_n3104), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__12_ ( .D(
        mem_stage_inst_dmem_n3105), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__13_ ( .D(
        mem_stage_inst_dmem_n3106), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__14_ ( .D(
        mem_stage_inst_dmem_n3107), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_158__15_ ( .D(
        mem_stage_inst_dmem_n3108), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_158__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__0_ ( .D(
        mem_stage_inst_dmem_n3157), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__1_ ( .D(
        mem_stage_inst_dmem_n3158), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__2_ ( .D(
        mem_stage_inst_dmem_n3159), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__3_ ( .D(
        mem_stage_inst_dmem_n3160), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__4_ ( .D(
        mem_stage_inst_dmem_n3161), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__5_ ( .D(
        mem_stage_inst_dmem_n3162), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__6_ ( .D(
        mem_stage_inst_dmem_n3163), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__7_ ( .D(
        mem_stage_inst_dmem_n3164), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__8_ ( .D(
        mem_stage_inst_dmem_n3165), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__9_ ( .D(
        mem_stage_inst_dmem_n3166), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__10_ ( .D(
        mem_stage_inst_dmem_n3167), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__11_ ( .D(
        mem_stage_inst_dmem_n3168), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__12_ ( .D(
        mem_stage_inst_dmem_n3169), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__13_ ( .D(
        mem_stage_inst_dmem_n3170), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__14_ ( .D(
        mem_stage_inst_dmem_n3171), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_162__15_ ( .D(
        mem_stage_inst_dmem_n3172), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_162__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__0_ ( .D(
        mem_stage_inst_dmem_n3221), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__1_ ( .D(
        mem_stage_inst_dmem_n3222), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__2_ ( .D(
        mem_stage_inst_dmem_n3223), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__3_ ( .D(
        mem_stage_inst_dmem_n3224), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__4_ ( .D(
        mem_stage_inst_dmem_n3225), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__5_ ( .D(
        mem_stage_inst_dmem_n3226), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__6_ ( .D(
        mem_stage_inst_dmem_n3227), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__7_ ( .D(
        mem_stage_inst_dmem_n3228), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__8_ ( .D(
        mem_stage_inst_dmem_n3229), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__9_ ( .D(
        mem_stage_inst_dmem_n3230), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__10_ ( .D(
        mem_stage_inst_dmem_n3231), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__11_ ( .D(
        mem_stage_inst_dmem_n3232), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__12_ ( .D(
        mem_stage_inst_dmem_n3233), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__13_ ( .D(
        mem_stage_inst_dmem_n3234), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__14_ ( .D(
        mem_stage_inst_dmem_n3235), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_166__15_ ( .D(
        mem_stage_inst_dmem_n3236), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_166__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__0_ ( .D(
        mem_stage_inst_dmem_n3285), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__1_ ( .D(
        mem_stage_inst_dmem_n3286), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__2_ ( .D(
        mem_stage_inst_dmem_n3287), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__3_ ( .D(
        mem_stage_inst_dmem_n3288), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__4_ ( .D(
        mem_stage_inst_dmem_n3289), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__5_ ( .D(
        mem_stage_inst_dmem_n3290), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__6_ ( .D(
        mem_stage_inst_dmem_n3291), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__7_ ( .D(
        mem_stage_inst_dmem_n3292), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__8_ ( .D(
        mem_stage_inst_dmem_n3293), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__9_ ( .D(
        mem_stage_inst_dmem_n3294), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__10_ ( .D(
        mem_stage_inst_dmem_n3295), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__11_ ( .D(
        mem_stage_inst_dmem_n3296), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__12_ ( .D(
        mem_stage_inst_dmem_n3297), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__13_ ( .D(
        mem_stage_inst_dmem_n3298), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__14_ ( .D(
        mem_stage_inst_dmem_n3299), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_170__15_ ( .D(
        mem_stage_inst_dmem_n3300), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_170__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__0_ ( .D(
        mem_stage_inst_dmem_n3349), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__1_ ( .D(
        mem_stage_inst_dmem_n3350), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__2_ ( .D(
        mem_stage_inst_dmem_n3351), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__3_ ( .D(
        mem_stage_inst_dmem_n3352), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__4_ ( .D(
        mem_stage_inst_dmem_n3353), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__5_ ( .D(
        mem_stage_inst_dmem_n3354), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__6_ ( .D(
        mem_stage_inst_dmem_n3355), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__7_ ( .D(
        mem_stage_inst_dmem_n3356), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__8_ ( .D(
        mem_stage_inst_dmem_n3357), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__9_ ( .D(
        mem_stage_inst_dmem_n3358), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__10_ ( .D(
        mem_stage_inst_dmem_n3359), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__11_ ( .D(
        mem_stage_inst_dmem_n3360), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__12_ ( .D(
        mem_stage_inst_dmem_n3361), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__13_ ( .D(
        mem_stage_inst_dmem_n3362), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__14_ ( .D(
        mem_stage_inst_dmem_n3363), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_174__15_ ( .D(
        mem_stage_inst_dmem_n3364), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_174__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__0_ ( .D(
        mem_stage_inst_dmem_n3413), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__1_ ( .D(
        mem_stage_inst_dmem_n3414), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__2_ ( .D(
        mem_stage_inst_dmem_n3415), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__3_ ( .D(
        mem_stage_inst_dmem_n3416), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__4_ ( .D(
        mem_stage_inst_dmem_n3417), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__5_ ( .D(
        mem_stage_inst_dmem_n3418), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__6_ ( .D(
        mem_stage_inst_dmem_n3419), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__7_ ( .D(
        mem_stage_inst_dmem_n3420), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__8_ ( .D(
        mem_stage_inst_dmem_n3421), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__9_ ( .D(
        mem_stage_inst_dmem_n3422), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__10_ ( .D(
        mem_stage_inst_dmem_n3423), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__11_ ( .D(
        mem_stage_inst_dmem_n3424), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__12_ ( .D(
        mem_stage_inst_dmem_n3425), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__13_ ( .D(
        mem_stage_inst_dmem_n3426), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__14_ ( .D(
        mem_stage_inst_dmem_n3427), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_178__15_ ( .D(
        mem_stage_inst_dmem_n3428), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_178__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__0_ ( .D(
        mem_stage_inst_dmem_n3477), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__1_ ( .D(
        mem_stage_inst_dmem_n3478), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__2_ ( .D(
        mem_stage_inst_dmem_n3479), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__3_ ( .D(
        mem_stage_inst_dmem_n3480), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__4_ ( .D(
        mem_stage_inst_dmem_n3481), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__5_ ( .D(
        mem_stage_inst_dmem_n3482), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__6_ ( .D(
        mem_stage_inst_dmem_n3483), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__7_ ( .D(
        mem_stage_inst_dmem_n3484), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__8_ ( .D(
        mem_stage_inst_dmem_n3485), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__9_ ( .D(
        mem_stage_inst_dmem_n3486), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__10_ ( .D(
        mem_stage_inst_dmem_n3487), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__11_ ( .D(
        mem_stage_inst_dmem_n3488), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__12_ ( .D(
        mem_stage_inst_dmem_n3489), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__13_ ( .D(
        mem_stage_inst_dmem_n3490), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__14_ ( .D(
        mem_stage_inst_dmem_n3491), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_182__15_ ( .D(
        mem_stage_inst_dmem_n3492), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_182__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__0_ ( .D(
        mem_stage_inst_dmem_n3541), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__1_ ( .D(
        mem_stage_inst_dmem_n3542), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__2_ ( .D(
        mem_stage_inst_dmem_n3543), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__3_ ( .D(
        mem_stage_inst_dmem_n3544), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__4_ ( .D(
        mem_stage_inst_dmem_n3545), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__5_ ( .D(
        mem_stage_inst_dmem_n3546), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__6_ ( .D(
        mem_stage_inst_dmem_n3547), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__7_ ( .D(
        mem_stage_inst_dmem_n3548), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__8_ ( .D(
        mem_stage_inst_dmem_n3549), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__9_ ( .D(
        mem_stage_inst_dmem_n3550), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__10_ ( .D(
        mem_stage_inst_dmem_n3551), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__11_ ( .D(
        mem_stage_inst_dmem_n3552), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__12_ ( .D(
        mem_stage_inst_dmem_n3553), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__13_ ( .D(
        mem_stage_inst_dmem_n3554), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__14_ ( .D(
        mem_stage_inst_dmem_n3555), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_186__15_ ( .D(
        mem_stage_inst_dmem_n3556), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_186__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__0_ ( .D(
        mem_stage_inst_dmem_n3605), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__1_ ( .D(
        mem_stage_inst_dmem_n3606), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__2_ ( .D(
        mem_stage_inst_dmem_n3607), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__3_ ( .D(
        mem_stage_inst_dmem_n3608), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__4_ ( .D(
        mem_stage_inst_dmem_n3609), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__5_ ( .D(
        mem_stage_inst_dmem_n3610), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__6_ ( .D(
        mem_stage_inst_dmem_n3611), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__7_ ( .D(
        mem_stage_inst_dmem_n3612), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__8_ ( .D(
        mem_stage_inst_dmem_n3613), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__9_ ( .D(
        mem_stage_inst_dmem_n3614), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__10_ ( .D(
        mem_stage_inst_dmem_n3615), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__11_ ( .D(
        mem_stage_inst_dmem_n3616), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__12_ ( .D(
        mem_stage_inst_dmem_n3617), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__13_ ( .D(
        mem_stage_inst_dmem_n3618), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__14_ ( .D(
        mem_stage_inst_dmem_n3619), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_190__15_ ( .D(
        mem_stage_inst_dmem_n3620), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_190__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__0_ ( .D(
        mem_stage_inst_dmem_n3669), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__1_ ( .D(
        mem_stage_inst_dmem_n3670), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__2_ ( .D(
        mem_stage_inst_dmem_n3671), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__3_ ( .D(
        mem_stage_inst_dmem_n3672), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__4_ ( .D(
        mem_stage_inst_dmem_n3673), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__5_ ( .D(
        mem_stage_inst_dmem_n3674), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__6_ ( .D(
        mem_stage_inst_dmem_n3675), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__7_ ( .D(
        mem_stage_inst_dmem_n3676), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__8_ ( .D(
        mem_stage_inst_dmem_n3677), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__9_ ( .D(
        mem_stage_inst_dmem_n3678), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__10_ ( .D(
        mem_stage_inst_dmem_n3679), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__11_ ( .D(
        mem_stage_inst_dmem_n3680), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__12_ ( .D(
        mem_stage_inst_dmem_n3681), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__13_ ( .D(
        mem_stage_inst_dmem_n3682), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__14_ ( .D(
        mem_stage_inst_dmem_n3683), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_194__15_ ( .D(
        mem_stage_inst_dmem_n3684), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_194__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__0_ ( .D(
        mem_stage_inst_dmem_n3733), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__1_ ( .D(
        mem_stage_inst_dmem_n3734), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__2_ ( .D(
        mem_stage_inst_dmem_n3735), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__3_ ( .D(
        mem_stage_inst_dmem_n3736), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__4_ ( .D(
        mem_stage_inst_dmem_n3737), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__5_ ( .D(
        mem_stage_inst_dmem_n3738), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__6_ ( .D(
        mem_stage_inst_dmem_n3739), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__7_ ( .D(
        mem_stage_inst_dmem_n3740), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__8_ ( .D(
        mem_stage_inst_dmem_n3741), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__9_ ( .D(
        mem_stage_inst_dmem_n3742), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__10_ ( .D(
        mem_stage_inst_dmem_n3743), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__11_ ( .D(
        mem_stage_inst_dmem_n3744), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__12_ ( .D(
        mem_stage_inst_dmem_n3745), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__13_ ( .D(
        mem_stage_inst_dmem_n3746), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__14_ ( .D(
        mem_stage_inst_dmem_n3747), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_198__15_ ( .D(
        mem_stage_inst_dmem_n3748), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_198__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__0_ ( .D(
        mem_stage_inst_dmem_n3797), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__1_ ( .D(
        mem_stage_inst_dmem_n3798), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__2_ ( .D(
        mem_stage_inst_dmem_n3799), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__3_ ( .D(
        mem_stage_inst_dmem_n3800), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__4_ ( .D(
        mem_stage_inst_dmem_n3801), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__5_ ( .D(
        mem_stage_inst_dmem_n3802), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__6_ ( .D(
        mem_stage_inst_dmem_n3803), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__7_ ( .D(
        mem_stage_inst_dmem_n3804), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__8_ ( .D(
        mem_stage_inst_dmem_n3805), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__9_ ( .D(
        mem_stage_inst_dmem_n3806), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__10_ ( .D(
        mem_stage_inst_dmem_n3807), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__11_ ( .D(
        mem_stage_inst_dmem_n3808), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__12_ ( .D(
        mem_stage_inst_dmem_n3809), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__13_ ( .D(
        mem_stage_inst_dmem_n3810), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__14_ ( .D(
        mem_stage_inst_dmem_n3811), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_202__15_ ( .D(
        mem_stage_inst_dmem_n3812), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_202__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__0_ ( .D(
        mem_stage_inst_dmem_n3861), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__1_ ( .D(
        mem_stage_inst_dmem_n3862), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__2_ ( .D(
        mem_stage_inst_dmem_n3863), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__3_ ( .D(
        mem_stage_inst_dmem_n3864), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__4_ ( .D(
        mem_stage_inst_dmem_n3865), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__5_ ( .D(
        mem_stage_inst_dmem_n3866), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__6_ ( .D(
        mem_stage_inst_dmem_n3867), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__7_ ( .D(
        mem_stage_inst_dmem_n3868), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__8_ ( .D(
        mem_stage_inst_dmem_n3869), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__9_ ( .D(
        mem_stage_inst_dmem_n3870), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__10_ ( .D(
        mem_stage_inst_dmem_n3871), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__11_ ( .D(
        mem_stage_inst_dmem_n3872), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__12_ ( .D(
        mem_stage_inst_dmem_n3873), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__13_ ( .D(
        mem_stage_inst_dmem_n3874), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__14_ ( .D(
        mem_stage_inst_dmem_n3875), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_206__15_ ( .D(
        mem_stage_inst_dmem_n3876), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_206__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__0_ ( .D(
        mem_stage_inst_dmem_n3925), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__1_ ( .D(
        mem_stage_inst_dmem_n3926), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__2_ ( .D(
        mem_stage_inst_dmem_n3927), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__3_ ( .D(
        mem_stage_inst_dmem_n3928), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__4_ ( .D(
        mem_stage_inst_dmem_n3929), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__5_ ( .D(
        mem_stage_inst_dmem_n3930), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__6_ ( .D(
        mem_stage_inst_dmem_n3931), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__7_ ( .D(
        mem_stage_inst_dmem_n3932), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__8_ ( .D(
        mem_stage_inst_dmem_n3933), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__9_ ( .D(
        mem_stage_inst_dmem_n3934), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__10_ ( .D(
        mem_stage_inst_dmem_n3935), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__11_ ( .D(
        mem_stage_inst_dmem_n3936), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__12_ ( .D(
        mem_stage_inst_dmem_n3937), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__13_ ( .D(
        mem_stage_inst_dmem_n3938), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__14_ ( .D(
        mem_stage_inst_dmem_n3939), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_210__15_ ( .D(
        mem_stage_inst_dmem_n3940), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_210__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__0_ ( .D(
        mem_stage_inst_dmem_n3989), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__1_ ( .D(
        mem_stage_inst_dmem_n3990), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__2_ ( .D(
        mem_stage_inst_dmem_n3991), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__3_ ( .D(
        mem_stage_inst_dmem_n3992), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__4_ ( .D(
        mem_stage_inst_dmem_n3993), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__5_ ( .D(
        mem_stage_inst_dmem_n3994), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__6_ ( .D(
        mem_stage_inst_dmem_n3995), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__7_ ( .D(
        mem_stage_inst_dmem_n3996), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__8_ ( .D(
        mem_stage_inst_dmem_n3997), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__9_ ( .D(
        mem_stage_inst_dmem_n3998), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__10_ ( .D(
        mem_stage_inst_dmem_n3999), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__11_ ( .D(
        mem_stage_inst_dmem_n4000), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__12_ ( .D(
        mem_stage_inst_dmem_n4001), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__13_ ( .D(
        mem_stage_inst_dmem_n4002), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__14_ ( .D(
        mem_stage_inst_dmem_n4003), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_214__15_ ( .D(
        mem_stage_inst_dmem_n4004), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_214__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__0_ ( .D(
        mem_stage_inst_dmem_n4053), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__1_ ( .D(
        mem_stage_inst_dmem_n4054), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__2_ ( .D(
        mem_stage_inst_dmem_n4055), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__3_ ( .D(
        mem_stage_inst_dmem_n4056), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__4_ ( .D(
        mem_stage_inst_dmem_n4057), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__5_ ( .D(
        mem_stage_inst_dmem_n4058), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__6_ ( .D(
        mem_stage_inst_dmem_n4059), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__7_ ( .D(
        mem_stage_inst_dmem_n4060), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__8_ ( .D(
        mem_stage_inst_dmem_n4061), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__9_ ( .D(
        mem_stage_inst_dmem_n4062), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__10_ ( .D(
        mem_stage_inst_dmem_n4063), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__11_ ( .D(
        mem_stage_inst_dmem_n4064), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__12_ ( .D(
        mem_stage_inst_dmem_n4065), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__13_ ( .D(
        mem_stage_inst_dmem_n4066), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__14_ ( .D(
        mem_stage_inst_dmem_n4067), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_218__15_ ( .D(
        mem_stage_inst_dmem_n4068), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_218__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__0_ ( .D(
        mem_stage_inst_dmem_n4117), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__1_ ( .D(
        mem_stage_inst_dmem_n4118), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__2_ ( .D(
        mem_stage_inst_dmem_n4119), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__3_ ( .D(
        mem_stage_inst_dmem_n4120), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__4_ ( .D(
        mem_stage_inst_dmem_n4121), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__5_ ( .D(
        mem_stage_inst_dmem_n4122), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__6_ ( .D(
        mem_stage_inst_dmem_n4123), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__7_ ( .D(
        mem_stage_inst_dmem_n4124), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__8_ ( .D(
        mem_stage_inst_dmem_n4125), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__9_ ( .D(
        mem_stage_inst_dmem_n4126), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__10_ ( .D(
        mem_stage_inst_dmem_n4127), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__11_ ( .D(
        mem_stage_inst_dmem_n4128), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__12_ ( .D(
        mem_stage_inst_dmem_n4129), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__13_ ( .D(
        mem_stage_inst_dmem_n4130), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__14_ ( .D(
        mem_stage_inst_dmem_n4131), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_222__15_ ( .D(
        mem_stage_inst_dmem_n4132), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_222__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__0_ ( .D(
        mem_stage_inst_dmem_n4181), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__1_ ( .D(
        mem_stage_inst_dmem_n4182), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__2_ ( .D(
        mem_stage_inst_dmem_n4183), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__3_ ( .D(
        mem_stage_inst_dmem_n4184), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__4_ ( .D(
        mem_stage_inst_dmem_n4185), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__5_ ( .D(
        mem_stage_inst_dmem_n4186), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__6_ ( .D(
        mem_stage_inst_dmem_n4187), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__7_ ( .D(
        mem_stage_inst_dmem_n4188), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__8_ ( .D(
        mem_stage_inst_dmem_n4189), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__9_ ( .D(
        mem_stage_inst_dmem_n4190), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__10_ ( .D(
        mem_stage_inst_dmem_n4191), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__11_ ( .D(
        mem_stage_inst_dmem_n4192), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__12_ ( .D(
        mem_stage_inst_dmem_n4193), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__13_ ( .D(
        mem_stage_inst_dmem_n4194), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__14_ ( .D(
        mem_stage_inst_dmem_n4195), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_226__15_ ( .D(
        mem_stage_inst_dmem_n4196), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_226__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__0_ ( .D(
        mem_stage_inst_dmem_n4245), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__1_ ( .D(
        mem_stage_inst_dmem_n4246), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__2_ ( .D(
        mem_stage_inst_dmem_n4247), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__3_ ( .D(
        mem_stage_inst_dmem_n4248), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__4_ ( .D(
        mem_stage_inst_dmem_n4249), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__5_ ( .D(
        mem_stage_inst_dmem_n4250), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__6_ ( .D(
        mem_stage_inst_dmem_n4251), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__7_ ( .D(
        mem_stage_inst_dmem_n4252), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__8_ ( .D(
        mem_stage_inst_dmem_n4253), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__9_ ( .D(
        mem_stage_inst_dmem_n4254), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__10_ ( .D(
        mem_stage_inst_dmem_n4255), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__11_ ( .D(
        mem_stage_inst_dmem_n4256), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__12_ ( .D(
        mem_stage_inst_dmem_n4257), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__13_ ( .D(
        mem_stage_inst_dmem_n4258), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__14_ ( .D(
        mem_stage_inst_dmem_n4259), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_230__15_ ( .D(
        mem_stage_inst_dmem_n4260), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_230__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__0_ ( .D(
        mem_stage_inst_dmem_n4309), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__1_ ( .D(
        mem_stage_inst_dmem_n4310), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__2_ ( .D(
        mem_stage_inst_dmem_n4311), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__3_ ( .D(
        mem_stage_inst_dmem_n4312), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__4_ ( .D(
        mem_stage_inst_dmem_n4313), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__5_ ( .D(
        mem_stage_inst_dmem_n4314), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__6_ ( .D(
        mem_stage_inst_dmem_n4315), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__7_ ( .D(
        mem_stage_inst_dmem_n4316), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__8_ ( .D(
        mem_stage_inst_dmem_n4317), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__9_ ( .D(
        mem_stage_inst_dmem_n4318), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__10_ ( .D(
        mem_stage_inst_dmem_n4319), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__11_ ( .D(
        mem_stage_inst_dmem_n4320), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__12_ ( .D(
        mem_stage_inst_dmem_n4321), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__13_ ( .D(
        mem_stage_inst_dmem_n4322), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__14_ ( .D(
        mem_stage_inst_dmem_n4323), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_234__15_ ( .D(
        mem_stage_inst_dmem_n4324), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_234__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__0_ ( .D(
        mem_stage_inst_dmem_n4373), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__1_ ( .D(
        mem_stage_inst_dmem_n4374), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__2_ ( .D(
        mem_stage_inst_dmem_n4375), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__3_ ( .D(
        mem_stage_inst_dmem_n4376), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__4_ ( .D(
        mem_stage_inst_dmem_n4377), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__5_ ( .D(
        mem_stage_inst_dmem_n4378), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__6_ ( .D(
        mem_stage_inst_dmem_n4379), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__7_ ( .D(
        mem_stage_inst_dmem_n4380), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__8_ ( .D(
        mem_stage_inst_dmem_n4381), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__9_ ( .D(
        mem_stage_inst_dmem_n4382), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__10_ ( .D(
        mem_stage_inst_dmem_n4383), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__11_ ( .D(
        mem_stage_inst_dmem_n4384), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__12_ ( .D(
        mem_stage_inst_dmem_n4385), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__13_ ( .D(
        mem_stage_inst_dmem_n4386), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__14_ ( .D(
        mem_stage_inst_dmem_n4387), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_238__15_ ( .D(
        mem_stage_inst_dmem_n4388), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_238__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__0_ ( .D(
        mem_stage_inst_dmem_n4437), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__1_ ( .D(
        mem_stage_inst_dmem_n4438), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__2_ ( .D(
        mem_stage_inst_dmem_n4439), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__3_ ( .D(
        mem_stage_inst_dmem_n4440), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__4_ ( .D(
        mem_stage_inst_dmem_n4441), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__5_ ( .D(
        mem_stage_inst_dmem_n4442), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__6_ ( .D(
        mem_stage_inst_dmem_n4443), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__7_ ( .D(
        mem_stage_inst_dmem_n4444), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__8_ ( .D(
        mem_stage_inst_dmem_n4445), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__9_ ( .D(
        mem_stage_inst_dmem_n4446), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__10_ ( .D(
        mem_stage_inst_dmem_n4447), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__11_ ( .D(
        mem_stage_inst_dmem_n4448), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__12_ ( .D(
        mem_stage_inst_dmem_n4449), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__13_ ( .D(
        mem_stage_inst_dmem_n4450), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__14_ ( .D(
        mem_stage_inst_dmem_n4451), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_242__15_ ( .D(
        mem_stage_inst_dmem_n4452), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_242__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__0_ ( .D(
        mem_stage_inst_dmem_n4501), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__1_ ( .D(
        mem_stage_inst_dmem_n4502), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__2_ ( .D(
        mem_stage_inst_dmem_n4503), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__3_ ( .D(
        mem_stage_inst_dmem_n4504), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__4_ ( .D(
        mem_stage_inst_dmem_n4505), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__5_ ( .D(
        mem_stage_inst_dmem_n4506), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__6_ ( .D(
        mem_stage_inst_dmem_n4507), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__7_ ( .D(
        mem_stage_inst_dmem_n4508), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__8_ ( .D(
        mem_stage_inst_dmem_n4509), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__9_ ( .D(
        mem_stage_inst_dmem_n4510), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__10_ ( .D(
        mem_stage_inst_dmem_n4511), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__11_ ( .D(
        mem_stage_inst_dmem_n4512), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__12_ ( .D(
        mem_stage_inst_dmem_n4513), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__13_ ( .D(
        mem_stage_inst_dmem_n4514), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__14_ ( .D(
        mem_stage_inst_dmem_n4515), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_246__15_ ( .D(
        mem_stage_inst_dmem_n4516), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_246__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__0_ ( .D(
        mem_stage_inst_dmem_n4565), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__1_ ( .D(
        mem_stage_inst_dmem_n4566), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__2_ ( .D(
        mem_stage_inst_dmem_n4567), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__3_ ( .D(
        mem_stage_inst_dmem_n4568), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__4_ ( .D(
        mem_stage_inst_dmem_n4569), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__5_ ( .D(
        mem_stage_inst_dmem_n4570), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__6_ ( .D(
        mem_stage_inst_dmem_n4571), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__7_ ( .D(
        mem_stage_inst_dmem_n4572), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__8_ ( .D(
        mem_stage_inst_dmem_n4573), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__9_ ( .D(
        mem_stage_inst_dmem_n4574), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__10_ ( .D(
        mem_stage_inst_dmem_n4575), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__11_ ( .D(
        mem_stage_inst_dmem_n4576), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__12_ ( .D(
        mem_stage_inst_dmem_n4577), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__13_ ( .D(
        mem_stage_inst_dmem_n4578), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__14_ ( .D(
        mem_stage_inst_dmem_n4579), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_250__15_ ( .D(
        mem_stage_inst_dmem_n4580), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_250__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__0_ ( .D(
        mem_stage_inst_dmem_n4629), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__1_ ( .D(
        mem_stage_inst_dmem_n4630), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__2_ ( .D(
        mem_stage_inst_dmem_n4631), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__3_ ( .D(
        mem_stage_inst_dmem_n4632), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__4_ ( .D(
        mem_stage_inst_dmem_n4633), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__5_ ( .D(
        mem_stage_inst_dmem_n4634), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__6_ ( .D(
        mem_stage_inst_dmem_n4635), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__7_ ( .D(
        mem_stage_inst_dmem_n4636), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__8_ ( .D(
        mem_stage_inst_dmem_n4637), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__9_ ( .D(
        mem_stage_inst_dmem_n4638), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__10_ ( .D(
        mem_stage_inst_dmem_n4639), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__11_ ( .D(
        mem_stage_inst_dmem_n4640), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__12_ ( .D(
        mem_stage_inst_dmem_n4641), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__13_ ( .D(
        mem_stage_inst_dmem_n4642), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__14_ ( .D(
        mem_stage_inst_dmem_n4643), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_254__15_ ( .D(
        mem_stage_inst_dmem_n4644), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_254__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__0_ ( .D(
        mem_stage_inst_dmem_n565), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__1_ ( .D(
        mem_stage_inst_dmem_n566), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__2_ ( .D(
        mem_stage_inst_dmem_n567), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__3_ ( .D(
        mem_stage_inst_dmem_n568), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__4_ ( .D(
        mem_stage_inst_dmem_n569), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__5_ ( .D(
        mem_stage_inst_dmem_n570), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__6_ ( .D(
        mem_stage_inst_dmem_n571), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__7_ ( .D(
        mem_stage_inst_dmem_n572), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__8_ ( .D(
        mem_stage_inst_dmem_n573), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__9_ ( .D(
        mem_stage_inst_dmem_n574), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__10_ ( .D(
        mem_stage_inst_dmem_n575), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__11_ ( .D(
        mem_stage_inst_dmem_n576), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__12_ ( .D(
        mem_stage_inst_dmem_n577), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__13_ ( .D(
        mem_stage_inst_dmem_n578), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__14_ ( .D(
        mem_stage_inst_dmem_n579), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_0__15_ ( .D(
        mem_stage_inst_dmem_n580), .CK(clk), .Q(mem_stage_inst_dmem_ram_0__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__0_ ( .D(
        mem_stage_inst_dmem_n629), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__1_ ( .D(
        mem_stage_inst_dmem_n630), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__2_ ( .D(
        mem_stage_inst_dmem_n631), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__3_ ( .D(
        mem_stage_inst_dmem_n632), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__4_ ( .D(
        mem_stage_inst_dmem_n633), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__5_ ( .D(
        mem_stage_inst_dmem_n634), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__6_ ( .D(
        mem_stage_inst_dmem_n635), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__7_ ( .D(
        mem_stage_inst_dmem_n636), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__8_ ( .D(
        mem_stage_inst_dmem_n637), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__9_ ( .D(
        mem_stage_inst_dmem_n638), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__10_ ( .D(
        mem_stage_inst_dmem_n639), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__11_ ( .D(
        mem_stage_inst_dmem_n640), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__12_ ( .D(
        mem_stage_inst_dmem_n641), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__13_ ( .D(
        mem_stage_inst_dmem_n642), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__14_ ( .D(
        mem_stage_inst_dmem_n643), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_4__15_ ( .D(
        mem_stage_inst_dmem_n644), .CK(clk), .Q(mem_stage_inst_dmem_ram_4__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__0_ ( .D(
        mem_stage_inst_dmem_n693), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__1_ ( .D(
        mem_stage_inst_dmem_n694), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__2_ ( .D(
        mem_stage_inst_dmem_n695), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__3_ ( .D(
        mem_stage_inst_dmem_n696), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__4_ ( .D(
        mem_stage_inst_dmem_n697), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__5_ ( .D(
        mem_stage_inst_dmem_n698), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__6_ ( .D(
        mem_stage_inst_dmem_n699), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__7_ ( .D(
        mem_stage_inst_dmem_n700), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__8_ ( .D(
        mem_stage_inst_dmem_n701), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__9_ ( .D(
        mem_stage_inst_dmem_n702), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__10_ ( .D(
        mem_stage_inst_dmem_n703), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__11_ ( .D(
        mem_stage_inst_dmem_n704), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__12_ ( .D(
        mem_stage_inst_dmem_n705), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__13_ ( .D(
        mem_stage_inst_dmem_n706), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__14_ ( .D(
        mem_stage_inst_dmem_n707), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_8__15_ ( .D(
        mem_stage_inst_dmem_n708), .CK(clk), .Q(mem_stage_inst_dmem_ram_8__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__0_ ( .D(
        mem_stage_inst_dmem_n757), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__1_ ( .D(
        mem_stage_inst_dmem_n758), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__2_ ( .D(
        mem_stage_inst_dmem_n759), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__3_ ( .D(
        mem_stage_inst_dmem_n760), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__4_ ( .D(
        mem_stage_inst_dmem_n761), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__5_ ( .D(
        mem_stage_inst_dmem_n762), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__6_ ( .D(
        mem_stage_inst_dmem_n763), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__7_ ( .D(
        mem_stage_inst_dmem_n764), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__8_ ( .D(
        mem_stage_inst_dmem_n765), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__9_ ( .D(
        mem_stage_inst_dmem_n766), .CK(clk), .Q(mem_stage_inst_dmem_ram_12__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__10_ ( .D(
        mem_stage_inst_dmem_n767), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_12__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__11_ ( .D(
        mem_stage_inst_dmem_n768), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_12__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__12_ ( .D(
        mem_stage_inst_dmem_n769), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_12__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__13_ ( .D(
        mem_stage_inst_dmem_n770), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_12__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__14_ ( .D(
        mem_stage_inst_dmem_n771), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_12__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_12__15_ ( .D(
        mem_stage_inst_dmem_n772), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_12__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__0_ ( .D(
        mem_stage_inst_dmem_n821), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__1_ ( .D(
        mem_stage_inst_dmem_n822), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__2_ ( .D(
        mem_stage_inst_dmem_n823), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__3_ ( .D(
        mem_stage_inst_dmem_n824), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__4_ ( .D(
        mem_stage_inst_dmem_n825), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__5_ ( .D(
        mem_stage_inst_dmem_n826), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__6_ ( .D(
        mem_stage_inst_dmem_n827), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__7_ ( .D(
        mem_stage_inst_dmem_n828), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__8_ ( .D(
        mem_stage_inst_dmem_n829), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__9_ ( .D(
        mem_stage_inst_dmem_n830), .CK(clk), .Q(mem_stage_inst_dmem_ram_16__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__10_ ( .D(
        mem_stage_inst_dmem_n831), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_16__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__11_ ( .D(
        mem_stage_inst_dmem_n832), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_16__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__12_ ( .D(
        mem_stage_inst_dmem_n833), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_16__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__13_ ( .D(
        mem_stage_inst_dmem_n834), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_16__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__14_ ( .D(
        mem_stage_inst_dmem_n835), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_16__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_16__15_ ( .D(
        mem_stage_inst_dmem_n836), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_16__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__0_ ( .D(
        mem_stage_inst_dmem_n885), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__1_ ( .D(
        mem_stage_inst_dmem_n886), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__2_ ( .D(
        mem_stage_inst_dmem_n887), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__3_ ( .D(
        mem_stage_inst_dmem_n888), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__4_ ( .D(
        mem_stage_inst_dmem_n889), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__5_ ( .D(
        mem_stage_inst_dmem_n890), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__6_ ( .D(
        mem_stage_inst_dmem_n891), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__7_ ( .D(
        mem_stage_inst_dmem_n892), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__8_ ( .D(
        mem_stage_inst_dmem_n893), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__9_ ( .D(
        mem_stage_inst_dmem_n894), .CK(clk), .Q(mem_stage_inst_dmem_ram_20__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__10_ ( .D(
        mem_stage_inst_dmem_n895), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_20__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__11_ ( .D(
        mem_stage_inst_dmem_n896), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_20__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__12_ ( .D(
        mem_stage_inst_dmem_n897), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_20__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__13_ ( .D(
        mem_stage_inst_dmem_n898), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_20__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__14_ ( .D(
        mem_stage_inst_dmem_n899), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_20__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_20__15_ ( .D(
        mem_stage_inst_dmem_n900), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_20__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__0_ ( .D(
        mem_stage_inst_dmem_n949), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__1_ ( .D(
        mem_stage_inst_dmem_n950), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__2_ ( .D(
        mem_stage_inst_dmem_n951), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__3_ ( .D(
        mem_stage_inst_dmem_n952), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__4_ ( .D(
        mem_stage_inst_dmem_n953), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__5_ ( .D(
        mem_stage_inst_dmem_n954), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__6_ ( .D(
        mem_stage_inst_dmem_n955), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__7_ ( .D(
        mem_stage_inst_dmem_n956), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__8_ ( .D(
        mem_stage_inst_dmem_n957), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__9_ ( .D(
        mem_stage_inst_dmem_n958), .CK(clk), .Q(mem_stage_inst_dmem_ram_24__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__10_ ( .D(
        mem_stage_inst_dmem_n959), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_24__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__11_ ( .D(
        mem_stage_inst_dmem_n960), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_24__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__12_ ( .D(
        mem_stage_inst_dmem_n961), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_24__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__13_ ( .D(
        mem_stage_inst_dmem_n962), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_24__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__14_ ( .D(
        mem_stage_inst_dmem_n963), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_24__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_24__15_ ( .D(
        mem_stage_inst_dmem_n964), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_24__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__0_ ( .D(
        mem_stage_inst_dmem_n1013), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__1_ ( .D(
        mem_stage_inst_dmem_n1014), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__2_ ( .D(
        mem_stage_inst_dmem_n1015), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__3_ ( .D(
        mem_stage_inst_dmem_n1016), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__4_ ( .D(
        mem_stage_inst_dmem_n1017), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__5_ ( .D(
        mem_stage_inst_dmem_n1018), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__6_ ( .D(
        mem_stage_inst_dmem_n1019), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__7_ ( .D(
        mem_stage_inst_dmem_n1020), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__8_ ( .D(
        mem_stage_inst_dmem_n1021), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__9_ ( .D(
        mem_stage_inst_dmem_n1022), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__10_ ( .D(
        mem_stage_inst_dmem_n1023), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__11_ ( .D(
        mem_stage_inst_dmem_n1024), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__12_ ( .D(
        mem_stage_inst_dmem_n1025), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__13_ ( .D(
        mem_stage_inst_dmem_n1026), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__14_ ( .D(
        mem_stage_inst_dmem_n1027), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_28__15_ ( .D(
        mem_stage_inst_dmem_n1028), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_28__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__0_ ( .D(
        mem_stage_inst_dmem_n1077), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__1_ ( .D(
        mem_stage_inst_dmem_n1078), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__2_ ( .D(
        mem_stage_inst_dmem_n1079), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__3_ ( .D(
        mem_stage_inst_dmem_n1080), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__4_ ( .D(
        mem_stage_inst_dmem_n1081), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__5_ ( .D(
        mem_stage_inst_dmem_n1082), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__6_ ( .D(
        mem_stage_inst_dmem_n1083), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__7_ ( .D(
        mem_stage_inst_dmem_n1084), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__8_ ( .D(
        mem_stage_inst_dmem_n1085), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__9_ ( .D(
        mem_stage_inst_dmem_n1086), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__10_ ( .D(
        mem_stage_inst_dmem_n1087), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__11_ ( .D(
        mem_stage_inst_dmem_n1088), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__12_ ( .D(
        mem_stage_inst_dmem_n1089), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__13_ ( .D(
        mem_stage_inst_dmem_n1090), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__14_ ( .D(
        mem_stage_inst_dmem_n1091), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_32__15_ ( .D(
        mem_stage_inst_dmem_n1092), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_32__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__0_ ( .D(
        mem_stage_inst_dmem_n1141), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__1_ ( .D(
        mem_stage_inst_dmem_n1142), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__2_ ( .D(
        mem_stage_inst_dmem_n1143), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__3_ ( .D(
        mem_stage_inst_dmem_n1144), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__4_ ( .D(
        mem_stage_inst_dmem_n1145), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__5_ ( .D(
        mem_stage_inst_dmem_n1146), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__6_ ( .D(
        mem_stage_inst_dmem_n1147), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__7_ ( .D(
        mem_stage_inst_dmem_n1148), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__8_ ( .D(
        mem_stage_inst_dmem_n1149), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__9_ ( .D(
        mem_stage_inst_dmem_n1150), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__10_ ( .D(
        mem_stage_inst_dmem_n1151), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__11_ ( .D(
        mem_stage_inst_dmem_n1152), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__12_ ( .D(
        mem_stage_inst_dmem_n1153), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__13_ ( .D(
        mem_stage_inst_dmem_n1154), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__14_ ( .D(
        mem_stage_inst_dmem_n1155), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_36__15_ ( .D(
        mem_stage_inst_dmem_n1156), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_36__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__0_ ( .D(
        mem_stage_inst_dmem_n1205), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__1_ ( .D(
        mem_stage_inst_dmem_n1206), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__2_ ( .D(
        mem_stage_inst_dmem_n1207), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__3_ ( .D(
        mem_stage_inst_dmem_n1208), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__4_ ( .D(
        mem_stage_inst_dmem_n1209), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__5_ ( .D(
        mem_stage_inst_dmem_n1210), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__6_ ( .D(
        mem_stage_inst_dmem_n1211), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__7_ ( .D(
        mem_stage_inst_dmem_n1212), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__8_ ( .D(
        mem_stage_inst_dmem_n1213), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__9_ ( .D(
        mem_stage_inst_dmem_n1214), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__10_ ( .D(
        mem_stage_inst_dmem_n1215), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__11_ ( .D(
        mem_stage_inst_dmem_n1216), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__12_ ( .D(
        mem_stage_inst_dmem_n1217), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__13_ ( .D(
        mem_stage_inst_dmem_n1218), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__14_ ( .D(
        mem_stage_inst_dmem_n1219), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_40__15_ ( .D(
        mem_stage_inst_dmem_n1220), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_40__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__0_ ( .D(
        mem_stage_inst_dmem_n1269), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__1_ ( .D(
        mem_stage_inst_dmem_n1270), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__2_ ( .D(
        mem_stage_inst_dmem_n1271), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__3_ ( .D(
        mem_stage_inst_dmem_n1272), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__4_ ( .D(
        mem_stage_inst_dmem_n1273), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__5_ ( .D(
        mem_stage_inst_dmem_n1274), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__6_ ( .D(
        mem_stage_inst_dmem_n1275), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__7_ ( .D(
        mem_stage_inst_dmem_n1276), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__8_ ( .D(
        mem_stage_inst_dmem_n1277), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__9_ ( .D(
        mem_stage_inst_dmem_n1278), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__10_ ( .D(
        mem_stage_inst_dmem_n1279), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__11_ ( .D(
        mem_stage_inst_dmem_n1280), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__12_ ( .D(
        mem_stage_inst_dmem_n1281), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__13_ ( .D(
        mem_stage_inst_dmem_n1282), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__14_ ( .D(
        mem_stage_inst_dmem_n1283), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_44__15_ ( .D(
        mem_stage_inst_dmem_n1284), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_44__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__0_ ( .D(
        mem_stage_inst_dmem_n1333), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__1_ ( .D(
        mem_stage_inst_dmem_n1334), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__2_ ( .D(
        mem_stage_inst_dmem_n1335), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__3_ ( .D(
        mem_stage_inst_dmem_n1336), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__4_ ( .D(
        mem_stage_inst_dmem_n1337), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__5_ ( .D(
        mem_stage_inst_dmem_n1338), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__6_ ( .D(
        mem_stage_inst_dmem_n1339), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__7_ ( .D(
        mem_stage_inst_dmem_n1340), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__8_ ( .D(
        mem_stage_inst_dmem_n1341), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__9_ ( .D(
        mem_stage_inst_dmem_n1342), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__10_ ( .D(
        mem_stage_inst_dmem_n1343), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__11_ ( .D(
        mem_stage_inst_dmem_n1344), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__12_ ( .D(
        mem_stage_inst_dmem_n1345), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__13_ ( .D(
        mem_stage_inst_dmem_n1346), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__14_ ( .D(
        mem_stage_inst_dmem_n1347), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_48__15_ ( .D(
        mem_stage_inst_dmem_n1348), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_48__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__0_ ( .D(
        mem_stage_inst_dmem_n1397), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__1_ ( .D(
        mem_stage_inst_dmem_n1398), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__2_ ( .D(
        mem_stage_inst_dmem_n1399), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__3_ ( .D(
        mem_stage_inst_dmem_n1400), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__4_ ( .D(
        mem_stage_inst_dmem_n1401), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__5_ ( .D(
        mem_stage_inst_dmem_n1402), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__6_ ( .D(
        mem_stage_inst_dmem_n1403), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__7_ ( .D(
        mem_stage_inst_dmem_n1404), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__8_ ( .D(
        mem_stage_inst_dmem_n1405), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__9_ ( .D(
        mem_stage_inst_dmem_n1406), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__10_ ( .D(
        mem_stage_inst_dmem_n1407), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__11_ ( .D(
        mem_stage_inst_dmem_n1408), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__12_ ( .D(
        mem_stage_inst_dmem_n1409), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__13_ ( .D(
        mem_stage_inst_dmem_n1410), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__14_ ( .D(
        mem_stage_inst_dmem_n1411), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_52__15_ ( .D(
        mem_stage_inst_dmem_n1412), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_52__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__0_ ( .D(
        mem_stage_inst_dmem_n1461), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__1_ ( .D(
        mem_stage_inst_dmem_n1462), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__2_ ( .D(
        mem_stage_inst_dmem_n1463), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__3_ ( .D(
        mem_stage_inst_dmem_n1464), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__4_ ( .D(
        mem_stage_inst_dmem_n1465), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__5_ ( .D(
        mem_stage_inst_dmem_n1466), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__6_ ( .D(
        mem_stage_inst_dmem_n1467), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__7_ ( .D(
        mem_stage_inst_dmem_n1468), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__8_ ( .D(
        mem_stage_inst_dmem_n1469), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__9_ ( .D(
        mem_stage_inst_dmem_n1470), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__10_ ( .D(
        mem_stage_inst_dmem_n1471), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__11_ ( .D(
        mem_stage_inst_dmem_n1472), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__12_ ( .D(
        mem_stage_inst_dmem_n1473), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__13_ ( .D(
        mem_stage_inst_dmem_n1474), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__14_ ( .D(
        mem_stage_inst_dmem_n1475), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_56__15_ ( .D(
        mem_stage_inst_dmem_n1476), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_56__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__0_ ( .D(
        mem_stage_inst_dmem_n1525), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__1_ ( .D(
        mem_stage_inst_dmem_n1526), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__2_ ( .D(
        mem_stage_inst_dmem_n1527), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__3_ ( .D(
        mem_stage_inst_dmem_n1528), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__4_ ( .D(
        mem_stage_inst_dmem_n1529), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__5_ ( .D(
        mem_stage_inst_dmem_n1530), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__6_ ( .D(
        mem_stage_inst_dmem_n1531), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__7_ ( .D(
        mem_stage_inst_dmem_n1532), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__8_ ( .D(
        mem_stage_inst_dmem_n1533), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__9_ ( .D(
        mem_stage_inst_dmem_n1534), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__10_ ( .D(
        mem_stage_inst_dmem_n1535), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__11_ ( .D(
        mem_stage_inst_dmem_n1536), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__12_ ( .D(
        mem_stage_inst_dmem_n1537), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__13_ ( .D(
        mem_stage_inst_dmem_n1538), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__14_ ( .D(
        mem_stage_inst_dmem_n1539), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_60__15_ ( .D(
        mem_stage_inst_dmem_n1540), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_60__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__0_ ( .D(
        mem_stage_inst_dmem_n1589), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__1_ ( .D(
        mem_stage_inst_dmem_n1590), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__2_ ( .D(
        mem_stage_inst_dmem_n1591), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__3_ ( .D(
        mem_stage_inst_dmem_n1592), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__4_ ( .D(
        mem_stage_inst_dmem_n1593), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__5_ ( .D(
        mem_stage_inst_dmem_n1594), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__6_ ( .D(
        mem_stage_inst_dmem_n1595), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__7_ ( .D(
        mem_stage_inst_dmem_n1596), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__8_ ( .D(
        mem_stage_inst_dmem_n1597), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__9_ ( .D(
        mem_stage_inst_dmem_n1598), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__10_ ( .D(
        mem_stage_inst_dmem_n1599), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__11_ ( .D(
        mem_stage_inst_dmem_n1600), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__12_ ( .D(
        mem_stage_inst_dmem_n1601), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__13_ ( .D(
        mem_stage_inst_dmem_n1602), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__14_ ( .D(
        mem_stage_inst_dmem_n1603), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_64__15_ ( .D(
        mem_stage_inst_dmem_n1604), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_64__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__0_ ( .D(
        mem_stage_inst_dmem_n1653), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__1_ ( .D(
        mem_stage_inst_dmem_n1654), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__2_ ( .D(
        mem_stage_inst_dmem_n1655), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__3_ ( .D(
        mem_stage_inst_dmem_n1656), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__4_ ( .D(
        mem_stage_inst_dmem_n1657), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__5_ ( .D(
        mem_stage_inst_dmem_n1658), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__6_ ( .D(
        mem_stage_inst_dmem_n1659), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__7_ ( .D(
        mem_stage_inst_dmem_n1660), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__8_ ( .D(
        mem_stage_inst_dmem_n1661), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__9_ ( .D(
        mem_stage_inst_dmem_n1662), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__10_ ( .D(
        mem_stage_inst_dmem_n1663), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__11_ ( .D(
        mem_stage_inst_dmem_n1664), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__12_ ( .D(
        mem_stage_inst_dmem_n1665), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__13_ ( .D(
        mem_stage_inst_dmem_n1666), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__14_ ( .D(
        mem_stage_inst_dmem_n1667), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_68__15_ ( .D(
        mem_stage_inst_dmem_n1668), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_68__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__0_ ( .D(
        mem_stage_inst_dmem_n1717), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__1_ ( .D(
        mem_stage_inst_dmem_n1718), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__2_ ( .D(
        mem_stage_inst_dmem_n1719), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__3_ ( .D(
        mem_stage_inst_dmem_n1720), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__4_ ( .D(
        mem_stage_inst_dmem_n1721), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__5_ ( .D(
        mem_stage_inst_dmem_n1722), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__6_ ( .D(
        mem_stage_inst_dmem_n1723), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__7_ ( .D(
        mem_stage_inst_dmem_n1724), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__8_ ( .D(
        mem_stage_inst_dmem_n1725), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__9_ ( .D(
        mem_stage_inst_dmem_n1726), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__10_ ( .D(
        mem_stage_inst_dmem_n1727), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__11_ ( .D(
        mem_stage_inst_dmem_n1728), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__12_ ( .D(
        mem_stage_inst_dmem_n1729), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__13_ ( .D(
        mem_stage_inst_dmem_n1730), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__14_ ( .D(
        mem_stage_inst_dmem_n1731), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_72__15_ ( .D(
        mem_stage_inst_dmem_n1732), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_72__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__0_ ( .D(
        mem_stage_inst_dmem_n1781), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__1_ ( .D(
        mem_stage_inst_dmem_n1782), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__2_ ( .D(
        mem_stage_inst_dmem_n1783), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__3_ ( .D(
        mem_stage_inst_dmem_n1784), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__4_ ( .D(
        mem_stage_inst_dmem_n1785), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__5_ ( .D(
        mem_stage_inst_dmem_n1786), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__6_ ( .D(
        mem_stage_inst_dmem_n1787), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__7_ ( .D(
        mem_stage_inst_dmem_n1788), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__8_ ( .D(
        mem_stage_inst_dmem_n1789), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__9_ ( .D(
        mem_stage_inst_dmem_n1790), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__10_ ( .D(
        mem_stage_inst_dmem_n1791), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__11_ ( .D(
        mem_stage_inst_dmem_n1792), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__12_ ( .D(
        mem_stage_inst_dmem_n1793), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__13_ ( .D(
        mem_stage_inst_dmem_n1794), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__14_ ( .D(
        mem_stage_inst_dmem_n1795), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_76__15_ ( .D(
        mem_stage_inst_dmem_n1796), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_76__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__0_ ( .D(
        mem_stage_inst_dmem_n1845), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__1_ ( .D(
        mem_stage_inst_dmem_n1846), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__2_ ( .D(
        mem_stage_inst_dmem_n1847), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__3_ ( .D(
        mem_stage_inst_dmem_n1848), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__4_ ( .D(
        mem_stage_inst_dmem_n1849), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__5_ ( .D(
        mem_stage_inst_dmem_n1850), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__6_ ( .D(
        mem_stage_inst_dmem_n1851), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__7_ ( .D(
        mem_stage_inst_dmem_n1852), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__8_ ( .D(
        mem_stage_inst_dmem_n1853), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__9_ ( .D(
        mem_stage_inst_dmem_n1854), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__10_ ( .D(
        mem_stage_inst_dmem_n1855), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__11_ ( .D(
        mem_stage_inst_dmem_n1856), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__12_ ( .D(
        mem_stage_inst_dmem_n1857), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__13_ ( .D(
        mem_stage_inst_dmem_n1858), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__14_ ( .D(
        mem_stage_inst_dmem_n1859), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_80__15_ ( .D(
        mem_stage_inst_dmem_n1860), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_80__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__0_ ( .D(
        mem_stage_inst_dmem_n1909), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__1_ ( .D(
        mem_stage_inst_dmem_n1910), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__2_ ( .D(
        mem_stage_inst_dmem_n1911), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__3_ ( .D(
        mem_stage_inst_dmem_n1912), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__4_ ( .D(
        mem_stage_inst_dmem_n1913), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__5_ ( .D(
        mem_stage_inst_dmem_n1914), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__6_ ( .D(
        mem_stage_inst_dmem_n1915), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__7_ ( .D(
        mem_stage_inst_dmem_n1916), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__8_ ( .D(
        mem_stage_inst_dmem_n1917), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__9_ ( .D(
        mem_stage_inst_dmem_n1918), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__10_ ( .D(
        mem_stage_inst_dmem_n1919), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__11_ ( .D(
        mem_stage_inst_dmem_n1920), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__12_ ( .D(
        mem_stage_inst_dmem_n1921), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__13_ ( .D(
        mem_stage_inst_dmem_n1922), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__14_ ( .D(
        mem_stage_inst_dmem_n1923), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_84__15_ ( .D(
        mem_stage_inst_dmem_n1924), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_84__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__0_ ( .D(
        mem_stage_inst_dmem_n1973), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__1_ ( .D(
        mem_stage_inst_dmem_n1974), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__2_ ( .D(
        mem_stage_inst_dmem_n1975), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__3_ ( .D(
        mem_stage_inst_dmem_n1976), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__4_ ( .D(
        mem_stage_inst_dmem_n1977), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__5_ ( .D(
        mem_stage_inst_dmem_n1978), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__6_ ( .D(
        mem_stage_inst_dmem_n1979), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__7_ ( .D(
        mem_stage_inst_dmem_n1980), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__8_ ( .D(
        mem_stage_inst_dmem_n1981), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__9_ ( .D(
        mem_stage_inst_dmem_n1982), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__10_ ( .D(
        mem_stage_inst_dmem_n1983), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__11_ ( .D(
        mem_stage_inst_dmem_n1984), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__12_ ( .D(
        mem_stage_inst_dmem_n1985), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__13_ ( .D(
        mem_stage_inst_dmem_n1986), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__14_ ( .D(
        mem_stage_inst_dmem_n1987), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_88__15_ ( .D(
        mem_stage_inst_dmem_n1988), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_88__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__0_ ( .D(
        mem_stage_inst_dmem_n2037), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__1_ ( .D(
        mem_stage_inst_dmem_n2038), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__2_ ( .D(
        mem_stage_inst_dmem_n2039), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__3_ ( .D(
        mem_stage_inst_dmem_n2040), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__4_ ( .D(
        mem_stage_inst_dmem_n2041), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__5_ ( .D(
        mem_stage_inst_dmem_n2042), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__6_ ( .D(
        mem_stage_inst_dmem_n2043), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__7_ ( .D(
        mem_stage_inst_dmem_n2044), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__8_ ( .D(
        mem_stage_inst_dmem_n2045), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__9_ ( .D(
        mem_stage_inst_dmem_n2046), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__10_ ( .D(
        mem_stage_inst_dmem_n2047), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__11_ ( .D(
        mem_stage_inst_dmem_n2048), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__12_ ( .D(
        mem_stage_inst_dmem_n2049), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__13_ ( .D(
        mem_stage_inst_dmem_n2050), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__14_ ( .D(
        mem_stage_inst_dmem_n2051), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_92__15_ ( .D(
        mem_stage_inst_dmem_n2052), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_92__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__0_ ( .D(
        mem_stage_inst_dmem_n2101), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__1_ ( .D(
        mem_stage_inst_dmem_n2102), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__2_ ( .D(
        mem_stage_inst_dmem_n2103), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__3_ ( .D(
        mem_stage_inst_dmem_n2104), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__4_ ( .D(
        mem_stage_inst_dmem_n2105), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__5_ ( .D(
        mem_stage_inst_dmem_n2106), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__6_ ( .D(
        mem_stage_inst_dmem_n2107), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__7_ ( .D(
        mem_stage_inst_dmem_n2108), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__8_ ( .D(
        mem_stage_inst_dmem_n2109), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__9_ ( .D(
        mem_stage_inst_dmem_n2110), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__10_ ( .D(
        mem_stage_inst_dmem_n2111), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__11_ ( .D(
        mem_stage_inst_dmem_n2112), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__12_ ( .D(
        mem_stage_inst_dmem_n2113), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__13_ ( .D(
        mem_stage_inst_dmem_n2114), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__14_ ( .D(
        mem_stage_inst_dmem_n2115), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_96__15_ ( .D(
        mem_stage_inst_dmem_n2116), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_96__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__0_ ( .D(
        mem_stage_inst_dmem_n2165), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__1_ ( .D(
        mem_stage_inst_dmem_n2166), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__2_ ( .D(
        mem_stage_inst_dmem_n2167), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__3_ ( .D(
        mem_stage_inst_dmem_n2168), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__4_ ( .D(
        mem_stage_inst_dmem_n2169), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__5_ ( .D(
        mem_stage_inst_dmem_n2170), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__6_ ( .D(
        mem_stage_inst_dmem_n2171), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__7_ ( .D(
        mem_stage_inst_dmem_n2172), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__8_ ( .D(
        mem_stage_inst_dmem_n2173), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__9_ ( .D(
        mem_stage_inst_dmem_n2174), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__10_ ( .D(
        mem_stage_inst_dmem_n2175), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__11_ ( .D(
        mem_stage_inst_dmem_n2176), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__12_ ( .D(
        mem_stage_inst_dmem_n2177), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__13_ ( .D(
        mem_stage_inst_dmem_n2178), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__14_ ( .D(
        mem_stage_inst_dmem_n2179), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_100__15_ ( .D(
        mem_stage_inst_dmem_n2180), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_100__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__0_ ( .D(
        mem_stage_inst_dmem_n2229), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__1_ ( .D(
        mem_stage_inst_dmem_n2230), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__2_ ( .D(
        mem_stage_inst_dmem_n2231), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__3_ ( .D(
        mem_stage_inst_dmem_n2232), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__4_ ( .D(
        mem_stage_inst_dmem_n2233), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__5_ ( .D(
        mem_stage_inst_dmem_n2234), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__6_ ( .D(
        mem_stage_inst_dmem_n2235), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__7_ ( .D(
        mem_stage_inst_dmem_n2236), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__8_ ( .D(
        mem_stage_inst_dmem_n2237), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__9_ ( .D(
        mem_stage_inst_dmem_n2238), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__10_ ( .D(
        mem_stage_inst_dmem_n2239), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__11_ ( .D(
        mem_stage_inst_dmem_n2240), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__12_ ( .D(
        mem_stage_inst_dmem_n2241), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__13_ ( .D(
        mem_stage_inst_dmem_n2242), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__14_ ( .D(
        mem_stage_inst_dmem_n2243), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_104__15_ ( .D(
        mem_stage_inst_dmem_n2244), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_104__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__0_ ( .D(
        mem_stage_inst_dmem_n2293), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__1_ ( .D(
        mem_stage_inst_dmem_n2294), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__2_ ( .D(
        mem_stage_inst_dmem_n2295), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__3_ ( .D(
        mem_stage_inst_dmem_n2296), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__4_ ( .D(
        mem_stage_inst_dmem_n2297), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__5_ ( .D(
        mem_stage_inst_dmem_n2298), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__6_ ( .D(
        mem_stage_inst_dmem_n2299), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__7_ ( .D(
        mem_stage_inst_dmem_n2300), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__8_ ( .D(
        mem_stage_inst_dmem_n2301), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__9_ ( .D(
        mem_stage_inst_dmem_n2302), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__10_ ( .D(
        mem_stage_inst_dmem_n2303), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__11_ ( .D(
        mem_stage_inst_dmem_n2304), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__12_ ( .D(
        mem_stage_inst_dmem_n2305), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__13_ ( .D(
        mem_stage_inst_dmem_n2306), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__14_ ( .D(
        mem_stage_inst_dmem_n2307), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_108__15_ ( .D(
        mem_stage_inst_dmem_n2308), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_108__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__0_ ( .D(
        mem_stage_inst_dmem_n2357), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__1_ ( .D(
        mem_stage_inst_dmem_n2358), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__2_ ( .D(
        mem_stage_inst_dmem_n2359), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__3_ ( .D(
        mem_stage_inst_dmem_n2360), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__4_ ( .D(
        mem_stage_inst_dmem_n2361), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__5_ ( .D(
        mem_stage_inst_dmem_n2362), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__6_ ( .D(
        mem_stage_inst_dmem_n2363), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__7_ ( .D(
        mem_stage_inst_dmem_n2364), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__8_ ( .D(
        mem_stage_inst_dmem_n2365), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__9_ ( .D(
        mem_stage_inst_dmem_n2366), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__10_ ( .D(
        mem_stage_inst_dmem_n2367), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__11_ ( .D(
        mem_stage_inst_dmem_n2368), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__12_ ( .D(
        mem_stage_inst_dmem_n2369), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__13_ ( .D(
        mem_stage_inst_dmem_n2370), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__14_ ( .D(
        mem_stage_inst_dmem_n2371), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_112__15_ ( .D(
        mem_stage_inst_dmem_n2372), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_112__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__0_ ( .D(
        mem_stage_inst_dmem_n2421), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__1_ ( .D(
        mem_stage_inst_dmem_n2422), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__2_ ( .D(
        mem_stage_inst_dmem_n2423), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__3_ ( .D(
        mem_stage_inst_dmem_n2424), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__4_ ( .D(
        mem_stage_inst_dmem_n2425), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__5_ ( .D(
        mem_stage_inst_dmem_n2426), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__6_ ( .D(
        mem_stage_inst_dmem_n2427), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__7_ ( .D(
        mem_stage_inst_dmem_n2428), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__8_ ( .D(
        mem_stage_inst_dmem_n2429), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__9_ ( .D(
        mem_stage_inst_dmem_n2430), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__10_ ( .D(
        mem_stage_inst_dmem_n2431), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__11_ ( .D(
        mem_stage_inst_dmem_n2432), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__12_ ( .D(
        mem_stage_inst_dmem_n2433), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__13_ ( .D(
        mem_stage_inst_dmem_n2434), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__14_ ( .D(
        mem_stage_inst_dmem_n2435), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_116__15_ ( .D(
        mem_stage_inst_dmem_n2436), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_116__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__0_ ( .D(
        mem_stage_inst_dmem_n2485), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__1_ ( .D(
        mem_stage_inst_dmem_n2486), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__2_ ( .D(
        mem_stage_inst_dmem_n2487), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__3_ ( .D(
        mem_stage_inst_dmem_n2488), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__4_ ( .D(
        mem_stage_inst_dmem_n2489), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__5_ ( .D(
        mem_stage_inst_dmem_n2490), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__6_ ( .D(
        mem_stage_inst_dmem_n2491), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__7_ ( .D(
        mem_stage_inst_dmem_n2492), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__8_ ( .D(
        mem_stage_inst_dmem_n2493), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__9_ ( .D(
        mem_stage_inst_dmem_n2494), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__10_ ( .D(
        mem_stage_inst_dmem_n2495), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__11_ ( .D(
        mem_stage_inst_dmem_n2496), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__12_ ( .D(
        mem_stage_inst_dmem_n2497), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__13_ ( .D(
        mem_stage_inst_dmem_n2498), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__14_ ( .D(
        mem_stage_inst_dmem_n2499), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_120__15_ ( .D(
        mem_stage_inst_dmem_n2500), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_120__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__0_ ( .D(
        mem_stage_inst_dmem_n2549), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__1_ ( .D(
        mem_stage_inst_dmem_n2550), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__2_ ( .D(
        mem_stage_inst_dmem_n2551), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__3_ ( .D(
        mem_stage_inst_dmem_n2552), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__4_ ( .D(
        mem_stage_inst_dmem_n2553), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__5_ ( .D(
        mem_stage_inst_dmem_n2554), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__6_ ( .D(
        mem_stage_inst_dmem_n2555), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__7_ ( .D(
        mem_stage_inst_dmem_n2556), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__8_ ( .D(
        mem_stage_inst_dmem_n2557), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__9_ ( .D(
        mem_stage_inst_dmem_n2558), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__10_ ( .D(
        mem_stage_inst_dmem_n2559), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__11_ ( .D(
        mem_stage_inst_dmem_n2560), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__12_ ( .D(
        mem_stage_inst_dmem_n2561), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__13_ ( .D(
        mem_stage_inst_dmem_n2562), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__14_ ( .D(
        mem_stage_inst_dmem_n2563), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_124__15_ ( .D(
        mem_stage_inst_dmem_n2564), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_124__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__0_ ( .D(
        mem_stage_inst_dmem_n2613), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__1_ ( .D(
        mem_stage_inst_dmem_n2614), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__2_ ( .D(
        mem_stage_inst_dmem_n2615), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__3_ ( .D(
        mem_stage_inst_dmem_n2616), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__4_ ( .D(
        mem_stage_inst_dmem_n2617), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__5_ ( .D(
        mem_stage_inst_dmem_n2618), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__6_ ( .D(
        mem_stage_inst_dmem_n2619), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__7_ ( .D(
        mem_stage_inst_dmem_n2620), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__8_ ( .D(
        mem_stage_inst_dmem_n2621), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__9_ ( .D(
        mem_stage_inst_dmem_n2622), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__10_ ( .D(
        mem_stage_inst_dmem_n2623), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__11_ ( .D(
        mem_stage_inst_dmem_n2624), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__12_ ( .D(
        mem_stage_inst_dmem_n2625), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__13_ ( .D(
        mem_stage_inst_dmem_n2626), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__14_ ( .D(
        mem_stage_inst_dmem_n2627), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_128__15_ ( .D(
        mem_stage_inst_dmem_n2628), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_128__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__0_ ( .D(
        mem_stage_inst_dmem_n2677), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__1_ ( .D(
        mem_stage_inst_dmem_n2678), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__2_ ( .D(
        mem_stage_inst_dmem_n2679), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__3_ ( .D(
        mem_stage_inst_dmem_n2680), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__4_ ( .D(
        mem_stage_inst_dmem_n2681), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__5_ ( .D(
        mem_stage_inst_dmem_n2682), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__6_ ( .D(
        mem_stage_inst_dmem_n2683), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__7_ ( .D(
        mem_stage_inst_dmem_n2684), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__8_ ( .D(
        mem_stage_inst_dmem_n2685), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__9_ ( .D(
        mem_stage_inst_dmem_n2686), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__10_ ( .D(
        mem_stage_inst_dmem_n2687), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__11_ ( .D(
        mem_stage_inst_dmem_n2688), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__12_ ( .D(
        mem_stage_inst_dmem_n2689), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__13_ ( .D(
        mem_stage_inst_dmem_n2690), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__14_ ( .D(
        mem_stage_inst_dmem_n2691), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_132__15_ ( .D(
        mem_stage_inst_dmem_n2692), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_132__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__0_ ( .D(
        mem_stage_inst_dmem_n2741), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__1_ ( .D(
        mem_stage_inst_dmem_n2742), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__2_ ( .D(
        mem_stage_inst_dmem_n2743), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__3_ ( .D(
        mem_stage_inst_dmem_n2744), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__4_ ( .D(
        mem_stage_inst_dmem_n2745), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__5_ ( .D(
        mem_stage_inst_dmem_n2746), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__6_ ( .D(
        mem_stage_inst_dmem_n2747), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__7_ ( .D(
        mem_stage_inst_dmem_n2748), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__8_ ( .D(
        mem_stage_inst_dmem_n2749), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__9_ ( .D(
        mem_stage_inst_dmem_n2750), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__10_ ( .D(
        mem_stage_inst_dmem_n2751), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__11_ ( .D(
        mem_stage_inst_dmem_n2752), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__12_ ( .D(
        mem_stage_inst_dmem_n2753), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__13_ ( .D(
        mem_stage_inst_dmem_n2754), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__14_ ( .D(
        mem_stage_inst_dmem_n2755), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_136__15_ ( .D(
        mem_stage_inst_dmem_n2756), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_136__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__0_ ( .D(
        mem_stage_inst_dmem_n2805), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__1_ ( .D(
        mem_stage_inst_dmem_n2806), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__2_ ( .D(
        mem_stage_inst_dmem_n2807), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__3_ ( .D(
        mem_stage_inst_dmem_n2808), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__4_ ( .D(
        mem_stage_inst_dmem_n2809), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__5_ ( .D(
        mem_stage_inst_dmem_n2810), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__6_ ( .D(
        mem_stage_inst_dmem_n2811), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__7_ ( .D(
        mem_stage_inst_dmem_n2812), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__8_ ( .D(
        mem_stage_inst_dmem_n2813), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__9_ ( .D(
        mem_stage_inst_dmem_n2814), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__10_ ( .D(
        mem_stage_inst_dmem_n2815), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__11_ ( .D(
        mem_stage_inst_dmem_n2816), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__12_ ( .D(
        mem_stage_inst_dmem_n2817), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__13_ ( .D(
        mem_stage_inst_dmem_n2818), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__14_ ( .D(
        mem_stage_inst_dmem_n2819), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_140__15_ ( .D(
        mem_stage_inst_dmem_n2820), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_140__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__0_ ( .D(
        mem_stage_inst_dmem_n2869), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__1_ ( .D(
        mem_stage_inst_dmem_n2870), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__2_ ( .D(
        mem_stage_inst_dmem_n2871), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__3_ ( .D(
        mem_stage_inst_dmem_n2872), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__4_ ( .D(
        mem_stage_inst_dmem_n2873), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__5_ ( .D(
        mem_stage_inst_dmem_n2874), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__6_ ( .D(
        mem_stage_inst_dmem_n2875), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__7_ ( .D(
        mem_stage_inst_dmem_n2876), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__8_ ( .D(
        mem_stage_inst_dmem_n2877), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__9_ ( .D(
        mem_stage_inst_dmem_n2878), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__10_ ( .D(
        mem_stage_inst_dmem_n2879), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__11_ ( .D(
        mem_stage_inst_dmem_n2880), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__12_ ( .D(
        mem_stage_inst_dmem_n2881), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__13_ ( .D(
        mem_stage_inst_dmem_n2882), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__14_ ( .D(
        mem_stage_inst_dmem_n2883), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_144__15_ ( .D(
        mem_stage_inst_dmem_n2884), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_144__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__0_ ( .D(
        mem_stage_inst_dmem_n2933), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__1_ ( .D(
        mem_stage_inst_dmem_n2934), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__2_ ( .D(
        mem_stage_inst_dmem_n2935), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__3_ ( .D(
        mem_stage_inst_dmem_n2936), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__4_ ( .D(
        mem_stage_inst_dmem_n2937), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__5_ ( .D(
        mem_stage_inst_dmem_n2938), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__6_ ( .D(
        mem_stage_inst_dmem_n2939), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__7_ ( .D(
        mem_stage_inst_dmem_n2940), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__8_ ( .D(
        mem_stage_inst_dmem_n2941), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__9_ ( .D(
        mem_stage_inst_dmem_n2942), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__10_ ( .D(
        mem_stage_inst_dmem_n2943), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__11_ ( .D(
        mem_stage_inst_dmem_n2944), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__12_ ( .D(
        mem_stage_inst_dmem_n2945), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__13_ ( .D(
        mem_stage_inst_dmem_n2946), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__14_ ( .D(
        mem_stage_inst_dmem_n2947), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_148__15_ ( .D(
        mem_stage_inst_dmem_n2948), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_148__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__0_ ( .D(
        mem_stage_inst_dmem_n2997), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__1_ ( .D(
        mem_stage_inst_dmem_n2998), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__2_ ( .D(
        mem_stage_inst_dmem_n2999), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__3_ ( .D(
        mem_stage_inst_dmem_n3000), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__4_ ( .D(
        mem_stage_inst_dmem_n3001), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__5_ ( .D(
        mem_stage_inst_dmem_n3002), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__6_ ( .D(
        mem_stage_inst_dmem_n3003), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__7_ ( .D(
        mem_stage_inst_dmem_n3004), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__8_ ( .D(
        mem_stage_inst_dmem_n3005), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__9_ ( .D(
        mem_stage_inst_dmem_n3006), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__10_ ( .D(
        mem_stage_inst_dmem_n3007), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__11_ ( .D(
        mem_stage_inst_dmem_n3008), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__12_ ( .D(
        mem_stage_inst_dmem_n3009), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__13_ ( .D(
        mem_stage_inst_dmem_n3010), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__14_ ( .D(
        mem_stage_inst_dmem_n3011), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_152__15_ ( .D(
        mem_stage_inst_dmem_n3012), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_152__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__0_ ( .D(
        mem_stage_inst_dmem_n3061), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__1_ ( .D(
        mem_stage_inst_dmem_n3062), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__2_ ( .D(
        mem_stage_inst_dmem_n3063), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__3_ ( .D(
        mem_stage_inst_dmem_n3064), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__4_ ( .D(
        mem_stage_inst_dmem_n3065), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__5_ ( .D(
        mem_stage_inst_dmem_n3066), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__6_ ( .D(
        mem_stage_inst_dmem_n3067), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__7_ ( .D(
        mem_stage_inst_dmem_n3068), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__8_ ( .D(
        mem_stage_inst_dmem_n3069), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__9_ ( .D(
        mem_stage_inst_dmem_n3070), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__10_ ( .D(
        mem_stage_inst_dmem_n3071), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__11_ ( .D(
        mem_stage_inst_dmem_n3072), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__12_ ( .D(
        mem_stage_inst_dmem_n3073), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__13_ ( .D(
        mem_stage_inst_dmem_n3074), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__14_ ( .D(
        mem_stage_inst_dmem_n3075), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_156__15_ ( .D(
        mem_stage_inst_dmem_n3076), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_156__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__0_ ( .D(
        mem_stage_inst_dmem_n3125), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__1_ ( .D(
        mem_stage_inst_dmem_n3126), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__2_ ( .D(
        mem_stage_inst_dmem_n3127), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__3_ ( .D(
        mem_stage_inst_dmem_n3128), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__4_ ( .D(
        mem_stage_inst_dmem_n3129), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__5_ ( .D(
        mem_stage_inst_dmem_n3130), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__6_ ( .D(
        mem_stage_inst_dmem_n3131), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__7_ ( .D(
        mem_stage_inst_dmem_n3132), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__8_ ( .D(
        mem_stage_inst_dmem_n3133), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__9_ ( .D(
        mem_stage_inst_dmem_n3134), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__10_ ( .D(
        mem_stage_inst_dmem_n3135), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__11_ ( .D(
        mem_stage_inst_dmem_n3136), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__12_ ( .D(
        mem_stage_inst_dmem_n3137), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__13_ ( .D(
        mem_stage_inst_dmem_n3138), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__14_ ( .D(
        mem_stage_inst_dmem_n3139), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_160__15_ ( .D(
        mem_stage_inst_dmem_n3140), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_160__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__0_ ( .D(
        mem_stage_inst_dmem_n3189), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__1_ ( .D(
        mem_stage_inst_dmem_n3190), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__2_ ( .D(
        mem_stage_inst_dmem_n3191), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__3_ ( .D(
        mem_stage_inst_dmem_n3192), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__4_ ( .D(
        mem_stage_inst_dmem_n3193), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__5_ ( .D(
        mem_stage_inst_dmem_n3194), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__6_ ( .D(
        mem_stage_inst_dmem_n3195), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__7_ ( .D(
        mem_stage_inst_dmem_n3196), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__8_ ( .D(
        mem_stage_inst_dmem_n3197), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__9_ ( .D(
        mem_stage_inst_dmem_n3198), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__10_ ( .D(
        mem_stage_inst_dmem_n3199), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__11_ ( .D(
        mem_stage_inst_dmem_n3200), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__12_ ( .D(
        mem_stage_inst_dmem_n3201), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__13_ ( .D(
        mem_stage_inst_dmem_n3202), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__14_ ( .D(
        mem_stage_inst_dmem_n3203), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_164__15_ ( .D(
        mem_stage_inst_dmem_n3204), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_164__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__0_ ( .D(
        mem_stage_inst_dmem_n3253), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__1_ ( .D(
        mem_stage_inst_dmem_n3254), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__2_ ( .D(
        mem_stage_inst_dmem_n3255), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__3_ ( .D(
        mem_stage_inst_dmem_n3256), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__4_ ( .D(
        mem_stage_inst_dmem_n3257), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__5_ ( .D(
        mem_stage_inst_dmem_n3258), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__6_ ( .D(
        mem_stage_inst_dmem_n3259), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__7_ ( .D(
        mem_stage_inst_dmem_n3260), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__8_ ( .D(
        mem_stage_inst_dmem_n3261), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__9_ ( .D(
        mem_stage_inst_dmem_n3262), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__10_ ( .D(
        mem_stage_inst_dmem_n3263), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__11_ ( .D(
        mem_stage_inst_dmem_n3264), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__12_ ( .D(
        mem_stage_inst_dmem_n3265), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__13_ ( .D(
        mem_stage_inst_dmem_n3266), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__14_ ( .D(
        mem_stage_inst_dmem_n3267), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_168__15_ ( .D(
        mem_stage_inst_dmem_n3268), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_168__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__0_ ( .D(
        mem_stage_inst_dmem_n3317), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__1_ ( .D(
        mem_stage_inst_dmem_n3318), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__2_ ( .D(
        mem_stage_inst_dmem_n3319), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__3_ ( .D(
        mem_stage_inst_dmem_n3320), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__4_ ( .D(
        mem_stage_inst_dmem_n3321), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__5_ ( .D(
        mem_stage_inst_dmem_n3322), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__6_ ( .D(
        mem_stage_inst_dmem_n3323), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__7_ ( .D(
        mem_stage_inst_dmem_n3324), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__8_ ( .D(
        mem_stage_inst_dmem_n3325), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__9_ ( .D(
        mem_stage_inst_dmem_n3326), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__10_ ( .D(
        mem_stage_inst_dmem_n3327), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__11_ ( .D(
        mem_stage_inst_dmem_n3328), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__12_ ( .D(
        mem_stage_inst_dmem_n3329), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__13_ ( .D(
        mem_stage_inst_dmem_n3330), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__14_ ( .D(
        mem_stage_inst_dmem_n3331), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_172__15_ ( .D(
        mem_stage_inst_dmem_n3332), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_172__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__0_ ( .D(
        mem_stage_inst_dmem_n3381), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__1_ ( .D(
        mem_stage_inst_dmem_n3382), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__2_ ( .D(
        mem_stage_inst_dmem_n3383), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__3_ ( .D(
        mem_stage_inst_dmem_n3384), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__4_ ( .D(
        mem_stage_inst_dmem_n3385), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__5_ ( .D(
        mem_stage_inst_dmem_n3386), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__6_ ( .D(
        mem_stage_inst_dmem_n3387), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__7_ ( .D(
        mem_stage_inst_dmem_n3388), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__8_ ( .D(
        mem_stage_inst_dmem_n3389), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__9_ ( .D(
        mem_stage_inst_dmem_n3390), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__10_ ( .D(
        mem_stage_inst_dmem_n3391), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__11_ ( .D(
        mem_stage_inst_dmem_n3392), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__12_ ( .D(
        mem_stage_inst_dmem_n3393), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__13_ ( .D(
        mem_stage_inst_dmem_n3394), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__14_ ( .D(
        mem_stage_inst_dmem_n3395), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_176__15_ ( .D(
        mem_stage_inst_dmem_n3396), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_176__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__0_ ( .D(
        mem_stage_inst_dmem_n3445), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__1_ ( .D(
        mem_stage_inst_dmem_n3446), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__2_ ( .D(
        mem_stage_inst_dmem_n3447), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__3_ ( .D(
        mem_stage_inst_dmem_n3448), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__4_ ( .D(
        mem_stage_inst_dmem_n3449), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__5_ ( .D(
        mem_stage_inst_dmem_n3450), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__6_ ( .D(
        mem_stage_inst_dmem_n3451), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__7_ ( .D(
        mem_stage_inst_dmem_n3452), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__8_ ( .D(
        mem_stage_inst_dmem_n3453), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__9_ ( .D(
        mem_stage_inst_dmem_n3454), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__10_ ( .D(
        mem_stage_inst_dmem_n3455), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__11_ ( .D(
        mem_stage_inst_dmem_n3456), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__12_ ( .D(
        mem_stage_inst_dmem_n3457), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__13_ ( .D(
        mem_stage_inst_dmem_n3458), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__14_ ( .D(
        mem_stage_inst_dmem_n3459), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_180__15_ ( .D(
        mem_stage_inst_dmem_n3460), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_180__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__0_ ( .D(
        mem_stage_inst_dmem_n3509), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__1_ ( .D(
        mem_stage_inst_dmem_n3510), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__2_ ( .D(
        mem_stage_inst_dmem_n3511), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__3_ ( .D(
        mem_stage_inst_dmem_n3512), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__4_ ( .D(
        mem_stage_inst_dmem_n3513), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__5_ ( .D(
        mem_stage_inst_dmem_n3514), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__6_ ( .D(
        mem_stage_inst_dmem_n3515), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__7_ ( .D(
        mem_stage_inst_dmem_n3516), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__8_ ( .D(
        mem_stage_inst_dmem_n3517), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__9_ ( .D(
        mem_stage_inst_dmem_n3518), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__10_ ( .D(
        mem_stage_inst_dmem_n3519), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__11_ ( .D(
        mem_stage_inst_dmem_n3520), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__12_ ( .D(
        mem_stage_inst_dmem_n3521), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__13_ ( .D(
        mem_stage_inst_dmem_n3522), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__14_ ( .D(
        mem_stage_inst_dmem_n3523), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_184__15_ ( .D(
        mem_stage_inst_dmem_n3524), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_184__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__0_ ( .D(
        mem_stage_inst_dmem_n3573), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__1_ ( .D(
        mem_stage_inst_dmem_n3574), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__2_ ( .D(
        mem_stage_inst_dmem_n3575), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__3_ ( .D(
        mem_stage_inst_dmem_n3576), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__4_ ( .D(
        mem_stage_inst_dmem_n3577), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__5_ ( .D(
        mem_stage_inst_dmem_n3578), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__6_ ( .D(
        mem_stage_inst_dmem_n3579), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__7_ ( .D(
        mem_stage_inst_dmem_n3580), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__8_ ( .D(
        mem_stage_inst_dmem_n3581), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__9_ ( .D(
        mem_stage_inst_dmem_n3582), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__10_ ( .D(
        mem_stage_inst_dmem_n3583), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__11_ ( .D(
        mem_stage_inst_dmem_n3584), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__12_ ( .D(
        mem_stage_inst_dmem_n3585), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__13_ ( .D(
        mem_stage_inst_dmem_n3586), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__14_ ( .D(
        mem_stage_inst_dmem_n3587), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_188__15_ ( .D(
        mem_stage_inst_dmem_n3588), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_188__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__0_ ( .D(
        mem_stage_inst_dmem_n3637), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__1_ ( .D(
        mem_stage_inst_dmem_n3638), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__2_ ( .D(
        mem_stage_inst_dmem_n3639), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__3_ ( .D(
        mem_stage_inst_dmem_n3640), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__4_ ( .D(
        mem_stage_inst_dmem_n3641), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__5_ ( .D(
        mem_stage_inst_dmem_n3642), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__6_ ( .D(
        mem_stage_inst_dmem_n3643), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__7_ ( .D(
        mem_stage_inst_dmem_n3644), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__8_ ( .D(
        mem_stage_inst_dmem_n3645), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__9_ ( .D(
        mem_stage_inst_dmem_n3646), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__10_ ( .D(
        mem_stage_inst_dmem_n3647), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__11_ ( .D(
        mem_stage_inst_dmem_n3648), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__12_ ( .D(
        mem_stage_inst_dmem_n3649), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__13_ ( .D(
        mem_stage_inst_dmem_n3650), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__14_ ( .D(
        mem_stage_inst_dmem_n3651), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_192__15_ ( .D(
        mem_stage_inst_dmem_n3652), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_192__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__0_ ( .D(
        mem_stage_inst_dmem_n3701), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__1_ ( .D(
        mem_stage_inst_dmem_n3702), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__2_ ( .D(
        mem_stage_inst_dmem_n3703), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__3_ ( .D(
        mem_stage_inst_dmem_n3704), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__4_ ( .D(
        mem_stage_inst_dmem_n3705), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__5_ ( .D(
        mem_stage_inst_dmem_n3706), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__6_ ( .D(
        mem_stage_inst_dmem_n3707), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__7_ ( .D(
        mem_stage_inst_dmem_n3708), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__8_ ( .D(
        mem_stage_inst_dmem_n3709), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__9_ ( .D(
        mem_stage_inst_dmem_n3710), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__10_ ( .D(
        mem_stage_inst_dmem_n3711), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__11_ ( .D(
        mem_stage_inst_dmem_n3712), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__12_ ( .D(
        mem_stage_inst_dmem_n3713), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__13_ ( .D(
        mem_stage_inst_dmem_n3714), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__14_ ( .D(
        mem_stage_inst_dmem_n3715), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_196__15_ ( .D(
        mem_stage_inst_dmem_n3716), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_196__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__0_ ( .D(
        mem_stage_inst_dmem_n3765), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__1_ ( .D(
        mem_stage_inst_dmem_n3766), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__2_ ( .D(
        mem_stage_inst_dmem_n3767), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__3_ ( .D(
        mem_stage_inst_dmem_n3768), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__4_ ( .D(
        mem_stage_inst_dmem_n3769), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__5_ ( .D(
        mem_stage_inst_dmem_n3770), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__6_ ( .D(
        mem_stage_inst_dmem_n3771), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__7_ ( .D(
        mem_stage_inst_dmem_n3772), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__8_ ( .D(
        mem_stage_inst_dmem_n3773), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__9_ ( .D(
        mem_stage_inst_dmem_n3774), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__10_ ( .D(
        mem_stage_inst_dmem_n3775), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__11_ ( .D(
        mem_stage_inst_dmem_n3776), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__12_ ( .D(
        mem_stage_inst_dmem_n3777), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__13_ ( .D(
        mem_stage_inst_dmem_n3778), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__14_ ( .D(
        mem_stage_inst_dmem_n3779), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_200__15_ ( .D(
        mem_stage_inst_dmem_n3780), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_200__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__0_ ( .D(
        mem_stage_inst_dmem_n3829), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__1_ ( .D(
        mem_stage_inst_dmem_n3830), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__2_ ( .D(
        mem_stage_inst_dmem_n3831), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__3_ ( .D(
        mem_stage_inst_dmem_n3832), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__4_ ( .D(
        mem_stage_inst_dmem_n3833), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__5_ ( .D(
        mem_stage_inst_dmem_n3834), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__6_ ( .D(
        mem_stage_inst_dmem_n3835), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__7_ ( .D(
        mem_stage_inst_dmem_n3836), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__8_ ( .D(
        mem_stage_inst_dmem_n3837), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__9_ ( .D(
        mem_stage_inst_dmem_n3838), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__10_ ( .D(
        mem_stage_inst_dmem_n3839), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__11_ ( .D(
        mem_stage_inst_dmem_n3840), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__12_ ( .D(
        mem_stage_inst_dmem_n3841), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__13_ ( .D(
        mem_stage_inst_dmem_n3842), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__14_ ( .D(
        mem_stage_inst_dmem_n3843), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_204__15_ ( .D(
        mem_stage_inst_dmem_n3844), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_204__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__0_ ( .D(
        mem_stage_inst_dmem_n3893), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__1_ ( .D(
        mem_stage_inst_dmem_n3894), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__2_ ( .D(
        mem_stage_inst_dmem_n3895), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__3_ ( .D(
        mem_stage_inst_dmem_n3896), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__4_ ( .D(
        mem_stage_inst_dmem_n3897), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__5_ ( .D(
        mem_stage_inst_dmem_n3898), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__6_ ( .D(
        mem_stage_inst_dmem_n3899), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__7_ ( .D(
        mem_stage_inst_dmem_n3900), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__8_ ( .D(
        mem_stage_inst_dmem_n3901), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__9_ ( .D(
        mem_stage_inst_dmem_n3902), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__10_ ( .D(
        mem_stage_inst_dmem_n3903), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__11_ ( .D(
        mem_stage_inst_dmem_n3904), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__12_ ( .D(
        mem_stage_inst_dmem_n3905), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__13_ ( .D(
        mem_stage_inst_dmem_n3906), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__14_ ( .D(
        mem_stage_inst_dmem_n3907), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_208__15_ ( .D(
        mem_stage_inst_dmem_n3908), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_208__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__0_ ( .D(
        mem_stage_inst_dmem_n3957), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__1_ ( .D(
        mem_stage_inst_dmem_n3958), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__2_ ( .D(
        mem_stage_inst_dmem_n3959), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__3_ ( .D(
        mem_stage_inst_dmem_n3960), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__4_ ( .D(
        mem_stage_inst_dmem_n3961), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__5_ ( .D(
        mem_stage_inst_dmem_n3962), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__6_ ( .D(
        mem_stage_inst_dmem_n3963), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__7_ ( .D(
        mem_stage_inst_dmem_n3964), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__8_ ( .D(
        mem_stage_inst_dmem_n3965), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__9_ ( .D(
        mem_stage_inst_dmem_n3966), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__10_ ( .D(
        mem_stage_inst_dmem_n3967), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__11_ ( .D(
        mem_stage_inst_dmem_n3968), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__12_ ( .D(
        mem_stage_inst_dmem_n3969), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__13_ ( .D(
        mem_stage_inst_dmem_n3970), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__14_ ( .D(
        mem_stage_inst_dmem_n3971), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_212__15_ ( .D(
        mem_stage_inst_dmem_n3972), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_212__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__0_ ( .D(
        mem_stage_inst_dmem_n4021), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__1_ ( .D(
        mem_stage_inst_dmem_n4022), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__2_ ( .D(
        mem_stage_inst_dmem_n4023), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__3_ ( .D(
        mem_stage_inst_dmem_n4024), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__4_ ( .D(
        mem_stage_inst_dmem_n4025), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__5_ ( .D(
        mem_stage_inst_dmem_n4026), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__6_ ( .D(
        mem_stage_inst_dmem_n4027), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__7_ ( .D(
        mem_stage_inst_dmem_n4028), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__8_ ( .D(
        mem_stage_inst_dmem_n4029), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__9_ ( .D(
        mem_stage_inst_dmem_n4030), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__10_ ( .D(
        mem_stage_inst_dmem_n4031), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__11_ ( .D(
        mem_stage_inst_dmem_n4032), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__12_ ( .D(
        mem_stage_inst_dmem_n4033), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__13_ ( .D(
        mem_stage_inst_dmem_n4034), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__14_ ( .D(
        mem_stage_inst_dmem_n4035), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_216__15_ ( .D(
        mem_stage_inst_dmem_n4036), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_216__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__0_ ( .D(
        mem_stage_inst_dmem_n4085), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__1_ ( .D(
        mem_stage_inst_dmem_n4086), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__2_ ( .D(
        mem_stage_inst_dmem_n4087), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__3_ ( .D(
        mem_stage_inst_dmem_n4088), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__4_ ( .D(
        mem_stage_inst_dmem_n4089), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__5_ ( .D(
        mem_stage_inst_dmem_n4090), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__6_ ( .D(
        mem_stage_inst_dmem_n4091), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__7_ ( .D(
        mem_stage_inst_dmem_n4092), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__8_ ( .D(
        mem_stage_inst_dmem_n4093), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__9_ ( .D(
        mem_stage_inst_dmem_n4094), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__10_ ( .D(
        mem_stage_inst_dmem_n4095), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__11_ ( .D(
        mem_stage_inst_dmem_n4096), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__12_ ( .D(
        mem_stage_inst_dmem_n4097), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__13_ ( .D(
        mem_stage_inst_dmem_n4098), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__14_ ( .D(
        mem_stage_inst_dmem_n4099), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_220__15_ ( .D(
        mem_stage_inst_dmem_n4100), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_220__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__0_ ( .D(
        mem_stage_inst_dmem_n4149), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__1_ ( .D(
        mem_stage_inst_dmem_n4150), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__2_ ( .D(
        mem_stage_inst_dmem_n4151), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__3_ ( .D(
        mem_stage_inst_dmem_n4152), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__4_ ( .D(
        mem_stage_inst_dmem_n4153), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__5_ ( .D(
        mem_stage_inst_dmem_n4154), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__6_ ( .D(
        mem_stage_inst_dmem_n4155), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__7_ ( .D(
        mem_stage_inst_dmem_n4156), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__8_ ( .D(
        mem_stage_inst_dmem_n4157), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__9_ ( .D(
        mem_stage_inst_dmem_n4158), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__10_ ( .D(
        mem_stage_inst_dmem_n4159), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__11_ ( .D(
        mem_stage_inst_dmem_n4160), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__12_ ( .D(
        mem_stage_inst_dmem_n4161), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__13_ ( .D(
        mem_stage_inst_dmem_n4162), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__14_ ( .D(
        mem_stage_inst_dmem_n4163), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_224__15_ ( .D(
        mem_stage_inst_dmem_n4164), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_224__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__0_ ( .D(
        mem_stage_inst_dmem_n4213), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__1_ ( .D(
        mem_stage_inst_dmem_n4214), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__2_ ( .D(
        mem_stage_inst_dmem_n4215), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__3_ ( .D(
        mem_stage_inst_dmem_n4216), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__4_ ( .D(
        mem_stage_inst_dmem_n4217), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__5_ ( .D(
        mem_stage_inst_dmem_n4218), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__6_ ( .D(
        mem_stage_inst_dmem_n4219), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__7_ ( .D(
        mem_stage_inst_dmem_n4220), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__8_ ( .D(
        mem_stage_inst_dmem_n4221), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__9_ ( .D(
        mem_stage_inst_dmem_n4222), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__10_ ( .D(
        mem_stage_inst_dmem_n4223), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__11_ ( .D(
        mem_stage_inst_dmem_n4224), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__12_ ( .D(
        mem_stage_inst_dmem_n4225), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__13_ ( .D(
        mem_stage_inst_dmem_n4226), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__14_ ( .D(
        mem_stage_inst_dmem_n4227), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_228__15_ ( .D(
        mem_stage_inst_dmem_n4228), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_228__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__0_ ( .D(
        mem_stage_inst_dmem_n4277), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__1_ ( .D(
        mem_stage_inst_dmem_n4278), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__2_ ( .D(
        mem_stage_inst_dmem_n4279), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__3_ ( .D(
        mem_stage_inst_dmem_n4280), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__4_ ( .D(
        mem_stage_inst_dmem_n4281), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__5_ ( .D(
        mem_stage_inst_dmem_n4282), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__6_ ( .D(
        mem_stage_inst_dmem_n4283), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__7_ ( .D(
        mem_stage_inst_dmem_n4284), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__8_ ( .D(
        mem_stage_inst_dmem_n4285), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__9_ ( .D(
        mem_stage_inst_dmem_n4286), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__10_ ( .D(
        mem_stage_inst_dmem_n4287), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__11_ ( .D(
        mem_stage_inst_dmem_n4288), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__12_ ( .D(
        mem_stage_inst_dmem_n4289), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__13_ ( .D(
        mem_stage_inst_dmem_n4290), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__14_ ( .D(
        mem_stage_inst_dmem_n4291), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_232__15_ ( .D(
        mem_stage_inst_dmem_n4292), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_232__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__0_ ( .D(
        mem_stage_inst_dmem_n4341), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__1_ ( .D(
        mem_stage_inst_dmem_n4342), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__2_ ( .D(
        mem_stage_inst_dmem_n4343), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__3_ ( .D(
        mem_stage_inst_dmem_n4344), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__4_ ( .D(
        mem_stage_inst_dmem_n4345), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__5_ ( .D(
        mem_stage_inst_dmem_n4346), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__6_ ( .D(
        mem_stage_inst_dmem_n4347), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__7_ ( .D(
        mem_stage_inst_dmem_n4348), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__8_ ( .D(
        mem_stage_inst_dmem_n4349), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__9_ ( .D(
        mem_stage_inst_dmem_n4350), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__10_ ( .D(
        mem_stage_inst_dmem_n4351), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__11_ ( .D(
        mem_stage_inst_dmem_n4352), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__12_ ( .D(
        mem_stage_inst_dmem_n4353), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__13_ ( .D(
        mem_stage_inst_dmem_n4354), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__14_ ( .D(
        mem_stage_inst_dmem_n4355), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_236__15_ ( .D(
        mem_stage_inst_dmem_n4356), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_236__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__0_ ( .D(
        mem_stage_inst_dmem_n4405), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__1_ ( .D(
        mem_stage_inst_dmem_n4406), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__2_ ( .D(
        mem_stage_inst_dmem_n4407), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__3_ ( .D(
        mem_stage_inst_dmem_n4408), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__4_ ( .D(
        mem_stage_inst_dmem_n4409), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__5_ ( .D(
        mem_stage_inst_dmem_n4410), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__6_ ( .D(
        mem_stage_inst_dmem_n4411), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__7_ ( .D(
        mem_stage_inst_dmem_n4412), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__8_ ( .D(
        mem_stage_inst_dmem_n4413), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__9_ ( .D(
        mem_stage_inst_dmem_n4414), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__10_ ( .D(
        mem_stage_inst_dmem_n4415), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__11_ ( .D(
        mem_stage_inst_dmem_n4416), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__12_ ( .D(
        mem_stage_inst_dmem_n4417), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__13_ ( .D(
        mem_stage_inst_dmem_n4418), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__14_ ( .D(
        mem_stage_inst_dmem_n4419), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_240__15_ ( .D(
        mem_stage_inst_dmem_n4420), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_240__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__0_ ( .D(
        mem_stage_inst_dmem_n4469), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__1_ ( .D(
        mem_stage_inst_dmem_n4470), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__2_ ( .D(
        mem_stage_inst_dmem_n4471), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__3_ ( .D(
        mem_stage_inst_dmem_n4472), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__4_ ( .D(
        mem_stage_inst_dmem_n4473), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__5_ ( .D(
        mem_stage_inst_dmem_n4474), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__6_ ( .D(
        mem_stage_inst_dmem_n4475), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__7_ ( .D(
        mem_stage_inst_dmem_n4476), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__8_ ( .D(
        mem_stage_inst_dmem_n4477), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__9_ ( .D(
        mem_stage_inst_dmem_n4478), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__10_ ( .D(
        mem_stage_inst_dmem_n4479), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__11_ ( .D(
        mem_stage_inst_dmem_n4480), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__12_ ( .D(
        mem_stage_inst_dmem_n4481), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__13_ ( .D(
        mem_stage_inst_dmem_n4482), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__14_ ( .D(
        mem_stage_inst_dmem_n4483), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_244__15_ ( .D(
        mem_stage_inst_dmem_n4484), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_244__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__0_ ( .D(
        mem_stage_inst_dmem_n4533), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__1_ ( .D(
        mem_stage_inst_dmem_n4534), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__2_ ( .D(
        mem_stage_inst_dmem_n4535), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__3_ ( .D(
        mem_stage_inst_dmem_n4536), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__4_ ( .D(
        mem_stage_inst_dmem_n4537), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__5_ ( .D(
        mem_stage_inst_dmem_n4538), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__6_ ( .D(
        mem_stage_inst_dmem_n4539), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__7_ ( .D(
        mem_stage_inst_dmem_n4540), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__8_ ( .D(
        mem_stage_inst_dmem_n4541), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__9_ ( .D(
        mem_stage_inst_dmem_n4542), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__10_ ( .D(
        mem_stage_inst_dmem_n4543), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__11_ ( .D(
        mem_stage_inst_dmem_n4544), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__12_ ( .D(
        mem_stage_inst_dmem_n4545), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__13_ ( .D(
        mem_stage_inst_dmem_n4546), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__14_ ( .D(
        mem_stage_inst_dmem_n4547), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_248__15_ ( .D(
        mem_stage_inst_dmem_n4548), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_248__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__0_ ( .D(
        mem_stage_inst_dmem_n4597), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__1_ ( .D(
        mem_stage_inst_dmem_n4598), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__2_ ( .D(
        mem_stage_inst_dmem_n4599), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__3_ ( .D(
        mem_stage_inst_dmem_n4600), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__4_ ( .D(
        mem_stage_inst_dmem_n4601), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__5_ ( .D(
        mem_stage_inst_dmem_n4602), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__6_ ( .D(
        mem_stage_inst_dmem_n4603), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__7_ ( .D(
        mem_stage_inst_dmem_n4604), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__8_ ( .D(
        mem_stage_inst_dmem_n4605), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__9_ ( .D(
        mem_stage_inst_dmem_n4606), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__10_ ( .D(
        mem_stage_inst_dmem_n4607), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__11_ ( .D(
        mem_stage_inst_dmem_n4608), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__12_ ( .D(
        mem_stage_inst_dmem_n4609), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__13_ ( .D(
        mem_stage_inst_dmem_n4610), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__14_ ( .D(
        mem_stage_inst_dmem_n4611), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_252__15_ ( .D(
        mem_stage_inst_dmem_n4612), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_252__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__0_ ( .D(
        mem_stage_inst_dmem_n581), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__1_ ( .D(
        mem_stage_inst_dmem_n582), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__2_ ( .D(
        mem_stage_inst_dmem_n583), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__3_ ( .D(
        mem_stage_inst_dmem_n584), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__4_ ( .D(
        mem_stage_inst_dmem_n585), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__5_ ( .D(
        mem_stage_inst_dmem_n586), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__6_ ( .D(
        mem_stage_inst_dmem_n587), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__7_ ( .D(
        mem_stage_inst_dmem_n588), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__8_ ( .D(
        mem_stage_inst_dmem_n589), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__9_ ( .D(
        mem_stage_inst_dmem_n590), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__10_ ( .D(
        mem_stage_inst_dmem_n591), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__11_ ( .D(
        mem_stage_inst_dmem_n592), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__12_ ( .D(
        mem_stage_inst_dmem_n593), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__13_ ( .D(
        mem_stage_inst_dmem_n594), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__14_ ( .D(
        mem_stage_inst_dmem_n595), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_1__15_ ( .D(
        mem_stage_inst_dmem_n596), .CK(clk), .Q(mem_stage_inst_dmem_ram_1__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__0_ ( .D(
        mem_stage_inst_dmem_n645), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__1_ ( .D(
        mem_stage_inst_dmem_n646), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__2_ ( .D(
        mem_stage_inst_dmem_n647), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__3_ ( .D(
        mem_stage_inst_dmem_n648), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__4_ ( .D(
        mem_stage_inst_dmem_n649), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__5_ ( .D(
        mem_stage_inst_dmem_n650), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__6_ ( .D(
        mem_stage_inst_dmem_n651), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__7_ ( .D(
        mem_stage_inst_dmem_n652), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__8_ ( .D(
        mem_stage_inst_dmem_n653), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__9_ ( .D(
        mem_stage_inst_dmem_n654), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__10_ ( .D(
        mem_stage_inst_dmem_n655), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__11_ ( .D(
        mem_stage_inst_dmem_n656), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__12_ ( .D(
        mem_stage_inst_dmem_n657), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__13_ ( .D(
        mem_stage_inst_dmem_n658), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__14_ ( .D(
        mem_stage_inst_dmem_n659), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_5__15_ ( .D(
        mem_stage_inst_dmem_n660), .CK(clk), .Q(mem_stage_inst_dmem_ram_5__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__0_ ( .D(
        mem_stage_inst_dmem_n709), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__1_ ( .D(
        mem_stage_inst_dmem_n710), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__2_ ( .D(
        mem_stage_inst_dmem_n711), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__3_ ( .D(
        mem_stage_inst_dmem_n712), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__4_ ( .D(
        mem_stage_inst_dmem_n713), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__5_ ( .D(
        mem_stage_inst_dmem_n714), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__6_ ( .D(
        mem_stage_inst_dmem_n715), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__7_ ( .D(
        mem_stage_inst_dmem_n716), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__8_ ( .D(
        mem_stage_inst_dmem_n717), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__9_ ( .D(
        mem_stage_inst_dmem_n718), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__10_ ( .D(
        mem_stage_inst_dmem_n719), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__11_ ( .D(
        mem_stage_inst_dmem_n720), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__12_ ( .D(
        mem_stage_inst_dmem_n721), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__13_ ( .D(
        mem_stage_inst_dmem_n722), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__14_ ( .D(
        mem_stage_inst_dmem_n723), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_9__15_ ( .D(
        mem_stage_inst_dmem_n724), .CK(clk), .Q(mem_stage_inst_dmem_ram_9__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__0_ ( .D(
        mem_stage_inst_dmem_n773), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__1_ ( .D(
        mem_stage_inst_dmem_n774), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__2_ ( .D(
        mem_stage_inst_dmem_n775), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__3_ ( .D(
        mem_stage_inst_dmem_n776), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__4_ ( .D(
        mem_stage_inst_dmem_n777), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__5_ ( .D(
        mem_stage_inst_dmem_n778), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__6_ ( .D(
        mem_stage_inst_dmem_n779), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__7_ ( .D(
        mem_stage_inst_dmem_n780), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__8_ ( .D(
        mem_stage_inst_dmem_n781), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__9_ ( .D(
        mem_stage_inst_dmem_n782), .CK(clk), .Q(mem_stage_inst_dmem_ram_13__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__10_ ( .D(
        mem_stage_inst_dmem_n783), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_13__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__11_ ( .D(
        mem_stage_inst_dmem_n784), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_13__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__12_ ( .D(
        mem_stage_inst_dmem_n785), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_13__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__13_ ( .D(
        mem_stage_inst_dmem_n786), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_13__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__14_ ( .D(
        mem_stage_inst_dmem_n787), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_13__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_13__15_ ( .D(
        mem_stage_inst_dmem_n788), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_13__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__0_ ( .D(
        mem_stage_inst_dmem_n837), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__1_ ( .D(
        mem_stage_inst_dmem_n838), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__2_ ( .D(
        mem_stage_inst_dmem_n839), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__3_ ( .D(
        mem_stage_inst_dmem_n840), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__4_ ( .D(
        mem_stage_inst_dmem_n841), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__5_ ( .D(
        mem_stage_inst_dmem_n842), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__6_ ( .D(
        mem_stage_inst_dmem_n843), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__7_ ( .D(
        mem_stage_inst_dmem_n844), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__8_ ( .D(
        mem_stage_inst_dmem_n845), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__9_ ( .D(
        mem_stage_inst_dmem_n846), .CK(clk), .Q(mem_stage_inst_dmem_ram_17__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__10_ ( .D(
        mem_stage_inst_dmem_n847), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_17__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__11_ ( .D(
        mem_stage_inst_dmem_n848), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_17__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__12_ ( .D(
        mem_stage_inst_dmem_n849), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_17__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__13_ ( .D(
        mem_stage_inst_dmem_n850), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_17__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__14_ ( .D(
        mem_stage_inst_dmem_n851), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_17__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_17__15_ ( .D(
        mem_stage_inst_dmem_n852), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_17__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__0_ ( .D(
        mem_stage_inst_dmem_n901), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__1_ ( .D(
        mem_stage_inst_dmem_n902), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__2_ ( .D(
        mem_stage_inst_dmem_n903), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__3_ ( .D(
        mem_stage_inst_dmem_n904), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__4_ ( .D(
        mem_stage_inst_dmem_n905), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__5_ ( .D(
        mem_stage_inst_dmem_n906), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__6_ ( .D(
        mem_stage_inst_dmem_n907), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__7_ ( .D(
        mem_stage_inst_dmem_n908), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__8_ ( .D(
        mem_stage_inst_dmem_n909), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__9_ ( .D(
        mem_stage_inst_dmem_n910), .CK(clk), .Q(mem_stage_inst_dmem_ram_21__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__10_ ( .D(
        mem_stage_inst_dmem_n911), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_21__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__11_ ( .D(
        mem_stage_inst_dmem_n912), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_21__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__12_ ( .D(
        mem_stage_inst_dmem_n913), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_21__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__13_ ( .D(
        mem_stage_inst_dmem_n914), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_21__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__14_ ( .D(
        mem_stage_inst_dmem_n915), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_21__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_21__15_ ( .D(
        mem_stage_inst_dmem_n916), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_21__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__0_ ( .D(
        mem_stage_inst_dmem_n965), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__1_ ( .D(
        mem_stage_inst_dmem_n966), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__2_ ( .D(
        mem_stage_inst_dmem_n967), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__3_ ( .D(
        mem_stage_inst_dmem_n968), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__4_ ( .D(
        mem_stage_inst_dmem_n969), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__5_ ( .D(
        mem_stage_inst_dmem_n970), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__6_ ( .D(
        mem_stage_inst_dmem_n971), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__7_ ( .D(
        mem_stage_inst_dmem_n972), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__8_ ( .D(
        mem_stage_inst_dmem_n973), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__9_ ( .D(
        mem_stage_inst_dmem_n974), .CK(clk), .Q(mem_stage_inst_dmem_ram_25__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__10_ ( .D(
        mem_stage_inst_dmem_n975), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_25__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__11_ ( .D(
        mem_stage_inst_dmem_n976), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_25__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__12_ ( .D(
        mem_stage_inst_dmem_n977), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_25__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__13_ ( .D(
        mem_stage_inst_dmem_n978), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_25__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__14_ ( .D(
        mem_stage_inst_dmem_n979), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_25__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_25__15_ ( .D(
        mem_stage_inst_dmem_n980), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_25__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__0_ ( .D(
        mem_stage_inst_dmem_n1029), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__1_ ( .D(
        mem_stage_inst_dmem_n1030), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__2_ ( .D(
        mem_stage_inst_dmem_n1031), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__3_ ( .D(
        mem_stage_inst_dmem_n1032), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__4_ ( .D(
        mem_stage_inst_dmem_n1033), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__5_ ( .D(
        mem_stage_inst_dmem_n1034), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__6_ ( .D(
        mem_stage_inst_dmem_n1035), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__7_ ( .D(
        mem_stage_inst_dmem_n1036), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__8_ ( .D(
        mem_stage_inst_dmem_n1037), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__9_ ( .D(
        mem_stage_inst_dmem_n1038), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__10_ ( .D(
        mem_stage_inst_dmem_n1039), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__11_ ( .D(
        mem_stage_inst_dmem_n1040), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__12_ ( .D(
        mem_stage_inst_dmem_n1041), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__13_ ( .D(
        mem_stage_inst_dmem_n1042), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__14_ ( .D(
        mem_stage_inst_dmem_n1043), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_29__15_ ( .D(
        mem_stage_inst_dmem_n1044), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_29__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__0_ ( .D(
        mem_stage_inst_dmem_n1093), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__1_ ( .D(
        mem_stage_inst_dmem_n1094), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__2_ ( .D(
        mem_stage_inst_dmem_n1095), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__3_ ( .D(
        mem_stage_inst_dmem_n1096), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__4_ ( .D(
        mem_stage_inst_dmem_n1097), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__5_ ( .D(
        mem_stage_inst_dmem_n1098), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__6_ ( .D(
        mem_stage_inst_dmem_n1099), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__7_ ( .D(
        mem_stage_inst_dmem_n1100), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__8_ ( .D(
        mem_stage_inst_dmem_n1101), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__9_ ( .D(
        mem_stage_inst_dmem_n1102), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__10_ ( .D(
        mem_stage_inst_dmem_n1103), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__11_ ( .D(
        mem_stage_inst_dmem_n1104), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__12_ ( .D(
        mem_stage_inst_dmem_n1105), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__13_ ( .D(
        mem_stage_inst_dmem_n1106), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__14_ ( .D(
        mem_stage_inst_dmem_n1107), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_33__15_ ( .D(
        mem_stage_inst_dmem_n1108), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_33__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__0_ ( .D(
        mem_stage_inst_dmem_n1157), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__1_ ( .D(
        mem_stage_inst_dmem_n1158), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__2_ ( .D(
        mem_stage_inst_dmem_n1159), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__3_ ( .D(
        mem_stage_inst_dmem_n1160), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__4_ ( .D(
        mem_stage_inst_dmem_n1161), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__5_ ( .D(
        mem_stage_inst_dmem_n1162), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__6_ ( .D(
        mem_stage_inst_dmem_n1163), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__7_ ( .D(
        mem_stage_inst_dmem_n1164), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__8_ ( .D(
        mem_stage_inst_dmem_n1165), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__9_ ( .D(
        mem_stage_inst_dmem_n1166), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__10_ ( .D(
        mem_stage_inst_dmem_n1167), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__11_ ( .D(
        mem_stage_inst_dmem_n1168), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__12_ ( .D(
        mem_stage_inst_dmem_n1169), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__13_ ( .D(
        mem_stage_inst_dmem_n1170), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__14_ ( .D(
        mem_stage_inst_dmem_n1171), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_37__15_ ( .D(
        mem_stage_inst_dmem_n1172), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_37__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__0_ ( .D(
        mem_stage_inst_dmem_n1221), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__1_ ( .D(
        mem_stage_inst_dmem_n1222), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__2_ ( .D(
        mem_stage_inst_dmem_n1223), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__3_ ( .D(
        mem_stage_inst_dmem_n1224), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__4_ ( .D(
        mem_stage_inst_dmem_n1225), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__5_ ( .D(
        mem_stage_inst_dmem_n1226), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__6_ ( .D(
        mem_stage_inst_dmem_n1227), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__7_ ( .D(
        mem_stage_inst_dmem_n1228), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__8_ ( .D(
        mem_stage_inst_dmem_n1229), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__9_ ( .D(
        mem_stage_inst_dmem_n1230), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__10_ ( .D(
        mem_stage_inst_dmem_n1231), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__11_ ( .D(
        mem_stage_inst_dmem_n1232), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__12_ ( .D(
        mem_stage_inst_dmem_n1233), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__13_ ( .D(
        mem_stage_inst_dmem_n1234), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__14_ ( .D(
        mem_stage_inst_dmem_n1235), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_41__15_ ( .D(
        mem_stage_inst_dmem_n1236), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_41__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__0_ ( .D(
        mem_stage_inst_dmem_n1285), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__1_ ( .D(
        mem_stage_inst_dmem_n1286), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__2_ ( .D(
        mem_stage_inst_dmem_n1287), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__3_ ( .D(
        mem_stage_inst_dmem_n1288), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__4_ ( .D(
        mem_stage_inst_dmem_n1289), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__5_ ( .D(
        mem_stage_inst_dmem_n1290), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__6_ ( .D(
        mem_stage_inst_dmem_n1291), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__7_ ( .D(
        mem_stage_inst_dmem_n1292), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__8_ ( .D(
        mem_stage_inst_dmem_n1293), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__9_ ( .D(
        mem_stage_inst_dmem_n1294), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__10_ ( .D(
        mem_stage_inst_dmem_n1295), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__11_ ( .D(
        mem_stage_inst_dmem_n1296), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__12_ ( .D(
        mem_stage_inst_dmem_n1297), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__13_ ( .D(
        mem_stage_inst_dmem_n1298), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__14_ ( .D(
        mem_stage_inst_dmem_n1299), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_45__15_ ( .D(
        mem_stage_inst_dmem_n1300), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_45__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__0_ ( .D(
        mem_stage_inst_dmem_n1349), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__1_ ( .D(
        mem_stage_inst_dmem_n1350), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__2_ ( .D(
        mem_stage_inst_dmem_n1351), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__3_ ( .D(
        mem_stage_inst_dmem_n1352), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__4_ ( .D(
        mem_stage_inst_dmem_n1353), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__5_ ( .D(
        mem_stage_inst_dmem_n1354), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__6_ ( .D(
        mem_stage_inst_dmem_n1355), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__7_ ( .D(
        mem_stage_inst_dmem_n1356), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__8_ ( .D(
        mem_stage_inst_dmem_n1357), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__9_ ( .D(
        mem_stage_inst_dmem_n1358), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__10_ ( .D(
        mem_stage_inst_dmem_n1359), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__11_ ( .D(
        mem_stage_inst_dmem_n1360), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__12_ ( .D(
        mem_stage_inst_dmem_n1361), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__13_ ( .D(
        mem_stage_inst_dmem_n1362), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__14_ ( .D(
        mem_stage_inst_dmem_n1363), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_49__15_ ( .D(
        mem_stage_inst_dmem_n1364), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_49__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__0_ ( .D(
        mem_stage_inst_dmem_n1413), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__1_ ( .D(
        mem_stage_inst_dmem_n1414), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__2_ ( .D(
        mem_stage_inst_dmem_n1415), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__3_ ( .D(
        mem_stage_inst_dmem_n1416), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__4_ ( .D(
        mem_stage_inst_dmem_n1417), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__5_ ( .D(
        mem_stage_inst_dmem_n1418), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__6_ ( .D(
        mem_stage_inst_dmem_n1419), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__7_ ( .D(
        mem_stage_inst_dmem_n1420), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__8_ ( .D(
        mem_stage_inst_dmem_n1421), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__9_ ( .D(
        mem_stage_inst_dmem_n1422), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__10_ ( .D(
        mem_stage_inst_dmem_n1423), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__11_ ( .D(
        mem_stage_inst_dmem_n1424), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__12_ ( .D(
        mem_stage_inst_dmem_n1425), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__13_ ( .D(
        mem_stage_inst_dmem_n1426), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__14_ ( .D(
        mem_stage_inst_dmem_n1427), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_53__15_ ( .D(
        mem_stage_inst_dmem_n1428), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_53__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__0_ ( .D(
        mem_stage_inst_dmem_n1477), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__1_ ( .D(
        mem_stage_inst_dmem_n1478), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__2_ ( .D(
        mem_stage_inst_dmem_n1479), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__3_ ( .D(
        mem_stage_inst_dmem_n1480), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__4_ ( .D(
        mem_stage_inst_dmem_n1481), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__5_ ( .D(
        mem_stage_inst_dmem_n1482), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__6_ ( .D(
        mem_stage_inst_dmem_n1483), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__7_ ( .D(
        mem_stage_inst_dmem_n1484), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__8_ ( .D(
        mem_stage_inst_dmem_n1485), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__9_ ( .D(
        mem_stage_inst_dmem_n1486), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__10_ ( .D(
        mem_stage_inst_dmem_n1487), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__11_ ( .D(
        mem_stage_inst_dmem_n1488), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__12_ ( .D(
        mem_stage_inst_dmem_n1489), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__13_ ( .D(
        mem_stage_inst_dmem_n1490), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__14_ ( .D(
        mem_stage_inst_dmem_n1491), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_57__15_ ( .D(
        mem_stage_inst_dmem_n1492), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_57__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__0_ ( .D(
        mem_stage_inst_dmem_n1541), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__1_ ( .D(
        mem_stage_inst_dmem_n1542), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__2_ ( .D(
        mem_stage_inst_dmem_n1543), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__3_ ( .D(
        mem_stage_inst_dmem_n1544), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__4_ ( .D(
        mem_stage_inst_dmem_n1545), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__5_ ( .D(
        mem_stage_inst_dmem_n1546), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__6_ ( .D(
        mem_stage_inst_dmem_n1547), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__7_ ( .D(
        mem_stage_inst_dmem_n1548), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__8_ ( .D(
        mem_stage_inst_dmem_n1549), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__9_ ( .D(
        mem_stage_inst_dmem_n1550), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__10_ ( .D(
        mem_stage_inst_dmem_n1551), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__11_ ( .D(
        mem_stage_inst_dmem_n1552), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__12_ ( .D(
        mem_stage_inst_dmem_n1553), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__13_ ( .D(
        mem_stage_inst_dmem_n1554), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__14_ ( .D(
        mem_stage_inst_dmem_n1555), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_61__15_ ( .D(
        mem_stage_inst_dmem_n1556), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_61__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__0_ ( .D(
        mem_stage_inst_dmem_n1605), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__1_ ( .D(
        mem_stage_inst_dmem_n1606), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__2_ ( .D(
        mem_stage_inst_dmem_n1607), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__3_ ( .D(
        mem_stage_inst_dmem_n1608), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__4_ ( .D(
        mem_stage_inst_dmem_n1609), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__5_ ( .D(
        mem_stage_inst_dmem_n1610), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__6_ ( .D(
        mem_stage_inst_dmem_n1611), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__7_ ( .D(
        mem_stage_inst_dmem_n1612), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__8_ ( .D(
        mem_stage_inst_dmem_n1613), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__9_ ( .D(
        mem_stage_inst_dmem_n1614), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__10_ ( .D(
        mem_stage_inst_dmem_n1615), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__11_ ( .D(
        mem_stage_inst_dmem_n1616), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__12_ ( .D(
        mem_stage_inst_dmem_n1617), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__13_ ( .D(
        mem_stage_inst_dmem_n1618), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__14_ ( .D(
        mem_stage_inst_dmem_n1619), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_65__15_ ( .D(
        mem_stage_inst_dmem_n1620), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_65__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__0_ ( .D(
        mem_stage_inst_dmem_n1669), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__1_ ( .D(
        mem_stage_inst_dmem_n1670), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__2_ ( .D(
        mem_stage_inst_dmem_n1671), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__3_ ( .D(
        mem_stage_inst_dmem_n1672), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__4_ ( .D(
        mem_stage_inst_dmem_n1673), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__5_ ( .D(
        mem_stage_inst_dmem_n1674), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__6_ ( .D(
        mem_stage_inst_dmem_n1675), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__7_ ( .D(
        mem_stage_inst_dmem_n1676), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__8_ ( .D(
        mem_stage_inst_dmem_n1677), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__9_ ( .D(
        mem_stage_inst_dmem_n1678), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__10_ ( .D(
        mem_stage_inst_dmem_n1679), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__11_ ( .D(
        mem_stage_inst_dmem_n1680), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__12_ ( .D(
        mem_stage_inst_dmem_n1681), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__13_ ( .D(
        mem_stage_inst_dmem_n1682), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__14_ ( .D(
        mem_stage_inst_dmem_n1683), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_69__15_ ( .D(
        mem_stage_inst_dmem_n1684), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_69__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__0_ ( .D(
        mem_stage_inst_dmem_n1733), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__1_ ( .D(
        mem_stage_inst_dmem_n1734), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__2_ ( .D(
        mem_stage_inst_dmem_n1735), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__3_ ( .D(
        mem_stage_inst_dmem_n1736), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__4_ ( .D(
        mem_stage_inst_dmem_n1737), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__5_ ( .D(
        mem_stage_inst_dmem_n1738), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__6_ ( .D(
        mem_stage_inst_dmem_n1739), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__7_ ( .D(
        mem_stage_inst_dmem_n1740), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__8_ ( .D(
        mem_stage_inst_dmem_n1741), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__9_ ( .D(
        mem_stage_inst_dmem_n1742), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__10_ ( .D(
        mem_stage_inst_dmem_n1743), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__11_ ( .D(
        mem_stage_inst_dmem_n1744), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__12_ ( .D(
        mem_stage_inst_dmem_n1745), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__13_ ( .D(
        mem_stage_inst_dmem_n1746), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__14_ ( .D(
        mem_stage_inst_dmem_n1747), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_73__15_ ( .D(
        mem_stage_inst_dmem_n1748), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_73__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__0_ ( .D(
        mem_stage_inst_dmem_n1797), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__1_ ( .D(
        mem_stage_inst_dmem_n1798), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__2_ ( .D(
        mem_stage_inst_dmem_n1799), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__3_ ( .D(
        mem_stage_inst_dmem_n1800), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__4_ ( .D(
        mem_stage_inst_dmem_n1801), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__5_ ( .D(
        mem_stage_inst_dmem_n1802), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__6_ ( .D(
        mem_stage_inst_dmem_n1803), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__7_ ( .D(
        mem_stage_inst_dmem_n1804), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__8_ ( .D(
        mem_stage_inst_dmem_n1805), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__9_ ( .D(
        mem_stage_inst_dmem_n1806), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__10_ ( .D(
        mem_stage_inst_dmem_n1807), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__11_ ( .D(
        mem_stage_inst_dmem_n1808), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__12_ ( .D(
        mem_stage_inst_dmem_n1809), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__13_ ( .D(
        mem_stage_inst_dmem_n1810), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__14_ ( .D(
        mem_stage_inst_dmem_n1811), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_77__15_ ( .D(
        mem_stage_inst_dmem_n1812), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_77__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__0_ ( .D(
        mem_stage_inst_dmem_n1861), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__1_ ( .D(
        mem_stage_inst_dmem_n1862), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__2_ ( .D(
        mem_stage_inst_dmem_n1863), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__3_ ( .D(
        mem_stage_inst_dmem_n1864), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__4_ ( .D(
        mem_stage_inst_dmem_n1865), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__5_ ( .D(
        mem_stage_inst_dmem_n1866), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__6_ ( .D(
        mem_stage_inst_dmem_n1867), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__7_ ( .D(
        mem_stage_inst_dmem_n1868), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__8_ ( .D(
        mem_stage_inst_dmem_n1869), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__9_ ( .D(
        mem_stage_inst_dmem_n1870), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__10_ ( .D(
        mem_stage_inst_dmem_n1871), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__11_ ( .D(
        mem_stage_inst_dmem_n1872), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__12_ ( .D(
        mem_stage_inst_dmem_n1873), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__13_ ( .D(
        mem_stage_inst_dmem_n1874), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__14_ ( .D(
        mem_stage_inst_dmem_n1875), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_81__15_ ( .D(
        mem_stage_inst_dmem_n1876), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_81__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__0_ ( .D(
        mem_stage_inst_dmem_n1925), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__1_ ( .D(
        mem_stage_inst_dmem_n1926), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__2_ ( .D(
        mem_stage_inst_dmem_n1927), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__3_ ( .D(
        mem_stage_inst_dmem_n1928), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__4_ ( .D(
        mem_stage_inst_dmem_n1929), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__5_ ( .D(
        mem_stage_inst_dmem_n1930), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__6_ ( .D(
        mem_stage_inst_dmem_n1931), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__7_ ( .D(
        mem_stage_inst_dmem_n1932), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__8_ ( .D(
        mem_stage_inst_dmem_n1933), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__9_ ( .D(
        mem_stage_inst_dmem_n1934), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__10_ ( .D(
        mem_stage_inst_dmem_n1935), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__11_ ( .D(
        mem_stage_inst_dmem_n1936), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__12_ ( .D(
        mem_stage_inst_dmem_n1937), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__13_ ( .D(
        mem_stage_inst_dmem_n1938), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__14_ ( .D(
        mem_stage_inst_dmem_n1939), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_85__15_ ( .D(
        mem_stage_inst_dmem_n1940), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_85__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__0_ ( .D(
        mem_stage_inst_dmem_n1989), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__1_ ( .D(
        mem_stage_inst_dmem_n1990), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__2_ ( .D(
        mem_stage_inst_dmem_n1991), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__3_ ( .D(
        mem_stage_inst_dmem_n1992), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__4_ ( .D(
        mem_stage_inst_dmem_n1993), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__5_ ( .D(
        mem_stage_inst_dmem_n1994), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__6_ ( .D(
        mem_stage_inst_dmem_n1995), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__7_ ( .D(
        mem_stage_inst_dmem_n1996), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__8_ ( .D(
        mem_stage_inst_dmem_n1997), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__9_ ( .D(
        mem_stage_inst_dmem_n1998), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__10_ ( .D(
        mem_stage_inst_dmem_n1999), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__11_ ( .D(
        mem_stage_inst_dmem_n2000), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__12_ ( .D(
        mem_stage_inst_dmem_n2001), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__13_ ( .D(
        mem_stage_inst_dmem_n2002), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__14_ ( .D(
        mem_stage_inst_dmem_n2003), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_89__15_ ( .D(
        mem_stage_inst_dmem_n2004), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_89__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__0_ ( .D(
        mem_stage_inst_dmem_n2053), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__1_ ( .D(
        mem_stage_inst_dmem_n2054), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__2_ ( .D(
        mem_stage_inst_dmem_n2055), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__3_ ( .D(
        mem_stage_inst_dmem_n2056), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__4_ ( .D(
        mem_stage_inst_dmem_n2057), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__5_ ( .D(
        mem_stage_inst_dmem_n2058), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__6_ ( .D(
        mem_stage_inst_dmem_n2059), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__7_ ( .D(
        mem_stage_inst_dmem_n2060), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__8_ ( .D(
        mem_stage_inst_dmem_n2061), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__9_ ( .D(
        mem_stage_inst_dmem_n2062), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__10_ ( .D(
        mem_stage_inst_dmem_n2063), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__11_ ( .D(
        mem_stage_inst_dmem_n2064), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__12_ ( .D(
        mem_stage_inst_dmem_n2065), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__13_ ( .D(
        mem_stage_inst_dmem_n2066), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__14_ ( .D(
        mem_stage_inst_dmem_n2067), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_93__15_ ( .D(
        mem_stage_inst_dmem_n2068), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_93__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__0_ ( .D(
        mem_stage_inst_dmem_n2117), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__1_ ( .D(
        mem_stage_inst_dmem_n2118), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__2_ ( .D(
        mem_stage_inst_dmem_n2119), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__3_ ( .D(
        mem_stage_inst_dmem_n2120), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__4_ ( .D(
        mem_stage_inst_dmem_n2121), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__5_ ( .D(
        mem_stage_inst_dmem_n2122), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__6_ ( .D(
        mem_stage_inst_dmem_n2123), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__7_ ( .D(
        mem_stage_inst_dmem_n2124), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__8_ ( .D(
        mem_stage_inst_dmem_n2125), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__9_ ( .D(
        mem_stage_inst_dmem_n2126), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__10_ ( .D(
        mem_stage_inst_dmem_n2127), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__11_ ( .D(
        mem_stage_inst_dmem_n2128), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__12_ ( .D(
        mem_stage_inst_dmem_n2129), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__13_ ( .D(
        mem_stage_inst_dmem_n2130), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__14_ ( .D(
        mem_stage_inst_dmem_n2131), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_97__15_ ( .D(
        mem_stage_inst_dmem_n2132), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_97__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__0_ ( .D(
        mem_stage_inst_dmem_n2181), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__1_ ( .D(
        mem_stage_inst_dmem_n2182), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__2_ ( .D(
        mem_stage_inst_dmem_n2183), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__3_ ( .D(
        mem_stage_inst_dmem_n2184), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__4_ ( .D(
        mem_stage_inst_dmem_n2185), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__5_ ( .D(
        mem_stage_inst_dmem_n2186), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__6_ ( .D(
        mem_stage_inst_dmem_n2187), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__7_ ( .D(
        mem_stage_inst_dmem_n2188), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__8_ ( .D(
        mem_stage_inst_dmem_n2189), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__9_ ( .D(
        mem_stage_inst_dmem_n2190), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__10_ ( .D(
        mem_stage_inst_dmem_n2191), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__11_ ( .D(
        mem_stage_inst_dmem_n2192), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__12_ ( .D(
        mem_stage_inst_dmem_n2193), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__13_ ( .D(
        mem_stage_inst_dmem_n2194), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__14_ ( .D(
        mem_stage_inst_dmem_n2195), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_101__15_ ( .D(
        mem_stage_inst_dmem_n2196), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_101__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__0_ ( .D(
        mem_stage_inst_dmem_n2245), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__1_ ( .D(
        mem_stage_inst_dmem_n2246), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__2_ ( .D(
        mem_stage_inst_dmem_n2247), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__3_ ( .D(
        mem_stage_inst_dmem_n2248), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__4_ ( .D(
        mem_stage_inst_dmem_n2249), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__5_ ( .D(
        mem_stage_inst_dmem_n2250), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__6_ ( .D(
        mem_stage_inst_dmem_n2251), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__7_ ( .D(
        mem_stage_inst_dmem_n2252), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__8_ ( .D(
        mem_stage_inst_dmem_n2253), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__9_ ( .D(
        mem_stage_inst_dmem_n2254), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__10_ ( .D(
        mem_stage_inst_dmem_n2255), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__11_ ( .D(
        mem_stage_inst_dmem_n2256), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__12_ ( .D(
        mem_stage_inst_dmem_n2257), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__13_ ( .D(
        mem_stage_inst_dmem_n2258), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__14_ ( .D(
        mem_stage_inst_dmem_n2259), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_105__15_ ( .D(
        mem_stage_inst_dmem_n2260), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_105__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__0_ ( .D(
        mem_stage_inst_dmem_n2309), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__1_ ( .D(
        mem_stage_inst_dmem_n2310), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__2_ ( .D(
        mem_stage_inst_dmem_n2311), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__3_ ( .D(
        mem_stage_inst_dmem_n2312), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__4_ ( .D(
        mem_stage_inst_dmem_n2313), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__5_ ( .D(
        mem_stage_inst_dmem_n2314), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__6_ ( .D(
        mem_stage_inst_dmem_n2315), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__7_ ( .D(
        mem_stage_inst_dmem_n2316), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__8_ ( .D(
        mem_stage_inst_dmem_n2317), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__9_ ( .D(
        mem_stage_inst_dmem_n2318), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__10_ ( .D(
        mem_stage_inst_dmem_n2319), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__11_ ( .D(
        mem_stage_inst_dmem_n2320), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__12_ ( .D(
        mem_stage_inst_dmem_n2321), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__13_ ( .D(
        mem_stage_inst_dmem_n2322), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__14_ ( .D(
        mem_stage_inst_dmem_n2323), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_109__15_ ( .D(
        mem_stage_inst_dmem_n2324), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_109__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__0_ ( .D(
        mem_stage_inst_dmem_n2373), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__1_ ( .D(
        mem_stage_inst_dmem_n2374), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__2_ ( .D(
        mem_stage_inst_dmem_n2375), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__3_ ( .D(
        mem_stage_inst_dmem_n2376), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__4_ ( .D(
        mem_stage_inst_dmem_n2377), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__5_ ( .D(
        mem_stage_inst_dmem_n2378), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__6_ ( .D(
        mem_stage_inst_dmem_n2379), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__7_ ( .D(
        mem_stage_inst_dmem_n2380), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__8_ ( .D(
        mem_stage_inst_dmem_n2381), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__9_ ( .D(
        mem_stage_inst_dmem_n2382), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__10_ ( .D(
        mem_stage_inst_dmem_n2383), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__11_ ( .D(
        mem_stage_inst_dmem_n2384), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__12_ ( .D(
        mem_stage_inst_dmem_n2385), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__13_ ( .D(
        mem_stage_inst_dmem_n2386), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__14_ ( .D(
        mem_stage_inst_dmem_n2387), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_113__15_ ( .D(
        mem_stage_inst_dmem_n2388), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_113__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__0_ ( .D(
        mem_stage_inst_dmem_n2437), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__1_ ( .D(
        mem_stage_inst_dmem_n2438), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__2_ ( .D(
        mem_stage_inst_dmem_n2439), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__3_ ( .D(
        mem_stage_inst_dmem_n2440), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__4_ ( .D(
        mem_stage_inst_dmem_n2441), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__5_ ( .D(
        mem_stage_inst_dmem_n2442), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__6_ ( .D(
        mem_stage_inst_dmem_n2443), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__7_ ( .D(
        mem_stage_inst_dmem_n2444), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__8_ ( .D(
        mem_stage_inst_dmem_n2445), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__9_ ( .D(
        mem_stage_inst_dmem_n2446), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__10_ ( .D(
        mem_stage_inst_dmem_n2447), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__11_ ( .D(
        mem_stage_inst_dmem_n2448), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__12_ ( .D(
        mem_stage_inst_dmem_n2449), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__13_ ( .D(
        mem_stage_inst_dmem_n2450), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__14_ ( .D(
        mem_stage_inst_dmem_n2451), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_117__15_ ( .D(
        mem_stage_inst_dmem_n2452), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_117__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__0_ ( .D(
        mem_stage_inst_dmem_n2501), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__1_ ( .D(
        mem_stage_inst_dmem_n2502), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__2_ ( .D(
        mem_stage_inst_dmem_n2503), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__3_ ( .D(
        mem_stage_inst_dmem_n2504), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__4_ ( .D(
        mem_stage_inst_dmem_n2505), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__5_ ( .D(
        mem_stage_inst_dmem_n2506), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__6_ ( .D(
        mem_stage_inst_dmem_n2507), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__7_ ( .D(
        mem_stage_inst_dmem_n2508), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__8_ ( .D(
        mem_stage_inst_dmem_n2509), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__9_ ( .D(
        mem_stage_inst_dmem_n2510), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__10_ ( .D(
        mem_stage_inst_dmem_n2511), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__11_ ( .D(
        mem_stage_inst_dmem_n2512), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__12_ ( .D(
        mem_stage_inst_dmem_n2513), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__13_ ( .D(
        mem_stage_inst_dmem_n2514), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__14_ ( .D(
        mem_stage_inst_dmem_n2515), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_121__15_ ( .D(
        mem_stage_inst_dmem_n2516), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_121__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__0_ ( .D(
        mem_stage_inst_dmem_n2565), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__1_ ( .D(
        mem_stage_inst_dmem_n2566), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__2_ ( .D(
        mem_stage_inst_dmem_n2567), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__3_ ( .D(
        mem_stage_inst_dmem_n2568), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__4_ ( .D(
        mem_stage_inst_dmem_n2569), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__5_ ( .D(
        mem_stage_inst_dmem_n2570), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__6_ ( .D(
        mem_stage_inst_dmem_n2571), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__7_ ( .D(
        mem_stage_inst_dmem_n2572), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__8_ ( .D(
        mem_stage_inst_dmem_n2573), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__9_ ( .D(
        mem_stage_inst_dmem_n2574), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__10_ ( .D(
        mem_stage_inst_dmem_n2575), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__11_ ( .D(
        mem_stage_inst_dmem_n2576), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__12_ ( .D(
        mem_stage_inst_dmem_n2577), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__13_ ( .D(
        mem_stage_inst_dmem_n2578), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__14_ ( .D(
        mem_stage_inst_dmem_n2579), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_125__15_ ( .D(
        mem_stage_inst_dmem_n2580), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_125__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__0_ ( .D(
        mem_stage_inst_dmem_n2629), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__1_ ( .D(
        mem_stage_inst_dmem_n2630), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__2_ ( .D(
        mem_stage_inst_dmem_n2631), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__3_ ( .D(
        mem_stage_inst_dmem_n2632), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__4_ ( .D(
        mem_stage_inst_dmem_n2633), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__5_ ( .D(
        mem_stage_inst_dmem_n2634), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__6_ ( .D(
        mem_stage_inst_dmem_n2635), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__7_ ( .D(
        mem_stage_inst_dmem_n2636), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__8_ ( .D(
        mem_stage_inst_dmem_n2637), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__9_ ( .D(
        mem_stage_inst_dmem_n2638), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__10_ ( .D(
        mem_stage_inst_dmem_n2639), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__11_ ( .D(
        mem_stage_inst_dmem_n2640), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__12_ ( .D(
        mem_stage_inst_dmem_n2641), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__13_ ( .D(
        mem_stage_inst_dmem_n2642), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__14_ ( .D(
        mem_stage_inst_dmem_n2643), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_129__15_ ( .D(
        mem_stage_inst_dmem_n2644), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_129__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__0_ ( .D(
        mem_stage_inst_dmem_n2693), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__1_ ( .D(
        mem_stage_inst_dmem_n2694), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__2_ ( .D(
        mem_stage_inst_dmem_n2695), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__3_ ( .D(
        mem_stage_inst_dmem_n2696), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__4_ ( .D(
        mem_stage_inst_dmem_n2697), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__5_ ( .D(
        mem_stage_inst_dmem_n2698), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__6_ ( .D(
        mem_stage_inst_dmem_n2699), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__7_ ( .D(
        mem_stage_inst_dmem_n2700), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__8_ ( .D(
        mem_stage_inst_dmem_n2701), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__9_ ( .D(
        mem_stage_inst_dmem_n2702), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__10_ ( .D(
        mem_stage_inst_dmem_n2703), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__11_ ( .D(
        mem_stage_inst_dmem_n2704), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__12_ ( .D(
        mem_stage_inst_dmem_n2705), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__13_ ( .D(
        mem_stage_inst_dmem_n2706), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__14_ ( .D(
        mem_stage_inst_dmem_n2707), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_133__15_ ( .D(
        mem_stage_inst_dmem_n2708), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_133__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__0_ ( .D(
        mem_stage_inst_dmem_n2757), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__1_ ( .D(
        mem_stage_inst_dmem_n2758), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__2_ ( .D(
        mem_stage_inst_dmem_n2759), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__3_ ( .D(
        mem_stage_inst_dmem_n2760), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__4_ ( .D(
        mem_stage_inst_dmem_n2761), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__5_ ( .D(
        mem_stage_inst_dmem_n2762), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__6_ ( .D(
        mem_stage_inst_dmem_n2763), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__7_ ( .D(
        mem_stage_inst_dmem_n2764), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__8_ ( .D(
        mem_stage_inst_dmem_n2765), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__9_ ( .D(
        mem_stage_inst_dmem_n2766), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__10_ ( .D(
        mem_stage_inst_dmem_n2767), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__11_ ( .D(
        mem_stage_inst_dmem_n2768), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__12_ ( .D(
        mem_stage_inst_dmem_n2769), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__13_ ( .D(
        mem_stage_inst_dmem_n2770), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__14_ ( .D(
        mem_stage_inst_dmem_n2771), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_137__15_ ( .D(
        mem_stage_inst_dmem_n2772), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_137__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__0_ ( .D(
        mem_stage_inst_dmem_n2821), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__1_ ( .D(
        mem_stage_inst_dmem_n2822), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__2_ ( .D(
        mem_stage_inst_dmem_n2823), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__3_ ( .D(
        mem_stage_inst_dmem_n2824), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__4_ ( .D(
        mem_stage_inst_dmem_n2825), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__5_ ( .D(
        mem_stage_inst_dmem_n2826), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__6_ ( .D(
        mem_stage_inst_dmem_n2827), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__7_ ( .D(
        mem_stage_inst_dmem_n2828), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__8_ ( .D(
        mem_stage_inst_dmem_n2829), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__9_ ( .D(
        mem_stage_inst_dmem_n2830), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__10_ ( .D(
        mem_stage_inst_dmem_n2831), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__11_ ( .D(
        mem_stage_inst_dmem_n2832), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__12_ ( .D(
        mem_stage_inst_dmem_n2833), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__13_ ( .D(
        mem_stage_inst_dmem_n2834), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__14_ ( .D(
        mem_stage_inst_dmem_n2835), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_141__15_ ( .D(
        mem_stage_inst_dmem_n2836), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_141__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__0_ ( .D(
        mem_stage_inst_dmem_n2885), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__1_ ( .D(
        mem_stage_inst_dmem_n2886), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__2_ ( .D(
        mem_stage_inst_dmem_n2887), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__3_ ( .D(
        mem_stage_inst_dmem_n2888), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__4_ ( .D(
        mem_stage_inst_dmem_n2889), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__5_ ( .D(
        mem_stage_inst_dmem_n2890), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__6_ ( .D(
        mem_stage_inst_dmem_n2891), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__7_ ( .D(
        mem_stage_inst_dmem_n2892), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__8_ ( .D(
        mem_stage_inst_dmem_n2893), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__9_ ( .D(
        mem_stage_inst_dmem_n2894), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__10_ ( .D(
        mem_stage_inst_dmem_n2895), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__11_ ( .D(
        mem_stage_inst_dmem_n2896), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__12_ ( .D(
        mem_stage_inst_dmem_n2897), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__13_ ( .D(
        mem_stage_inst_dmem_n2898), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__14_ ( .D(
        mem_stage_inst_dmem_n2899), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_145__15_ ( .D(
        mem_stage_inst_dmem_n2900), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_145__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__0_ ( .D(
        mem_stage_inst_dmem_n2949), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__1_ ( .D(
        mem_stage_inst_dmem_n2950), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__2_ ( .D(
        mem_stage_inst_dmem_n2951), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__3_ ( .D(
        mem_stage_inst_dmem_n2952), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__4_ ( .D(
        mem_stage_inst_dmem_n2953), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__5_ ( .D(
        mem_stage_inst_dmem_n2954), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__6_ ( .D(
        mem_stage_inst_dmem_n2955), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__7_ ( .D(
        mem_stage_inst_dmem_n2956), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__8_ ( .D(
        mem_stage_inst_dmem_n2957), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__9_ ( .D(
        mem_stage_inst_dmem_n2958), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__10_ ( .D(
        mem_stage_inst_dmem_n2959), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__11_ ( .D(
        mem_stage_inst_dmem_n2960), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__12_ ( .D(
        mem_stage_inst_dmem_n2961), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__13_ ( .D(
        mem_stage_inst_dmem_n2962), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__14_ ( .D(
        mem_stage_inst_dmem_n2963), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_149__15_ ( .D(
        mem_stage_inst_dmem_n2964), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_149__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__0_ ( .D(
        mem_stage_inst_dmem_n3013), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__1_ ( .D(
        mem_stage_inst_dmem_n3014), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__2_ ( .D(
        mem_stage_inst_dmem_n3015), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__3_ ( .D(
        mem_stage_inst_dmem_n3016), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__4_ ( .D(
        mem_stage_inst_dmem_n3017), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__5_ ( .D(
        mem_stage_inst_dmem_n3018), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__6_ ( .D(
        mem_stage_inst_dmem_n3019), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__7_ ( .D(
        mem_stage_inst_dmem_n3020), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__8_ ( .D(
        mem_stage_inst_dmem_n3021), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__9_ ( .D(
        mem_stage_inst_dmem_n3022), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__10_ ( .D(
        mem_stage_inst_dmem_n3023), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__11_ ( .D(
        mem_stage_inst_dmem_n3024), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__12_ ( .D(
        mem_stage_inst_dmem_n3025), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__13_ ( .D(
        mem_stage_inst_dmem_n3026), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__14_ ( .D(
        mem_stage_inst_dmem_n3027), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_153__15_ ( .D(
        mem_stage_inst_dmem_n3028), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_153__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__0_ ( .D(
        mem_stage_inst_dmem_n3077), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__1_ ( .D(
        mem_stage_inst_dmem_n3078), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__2_ ( .D(
        mem_stage_inst_dmem_n3079), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__3_ ( .D(
        mem_stage_inst_dmem_n3080), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__4_ ( .D(
        mem_stage_inst_dmem_n3081), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__5_ ( .D(
        mem_stage_inst_dmem_n3082), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__6_ ( .D(
        mem_stage_inst_dmem_n3083), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__7_ ( .D(
        mem_stage_inst_dmem_n3084), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__8_ ( .D(
        mem_stage_inst_dmem_n3085), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__9_ ( .D(
        mem_stage_inst_dmem_n3086), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__10_ ( .D(
        mem_stage_inst_dmem_n3087), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__11_ ( .D(
        mem_stage_inst_dmem_n3088), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__12_ ( .D(
        mem_stage_inst_dmem_n3089), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__13_ ( .D(
        mem_stage_inst_dmem_n3090), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__14_ ( .D(
        mem_stage_inst_dmem_n3091), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_157__15_ ( .D(
        mem_stage_inst_dmem_n3092), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_157__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__0_ ( .D(
        mem_stage_inst_dmem_n3141), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__1_ ( .D(
        mem_stage_inst_dmem_n3142), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__2_ ( .D(
        mem_stage_inst_dmem_n3143), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__3_ ( .D(
        mem_stage_inst_dmem_n3144), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__4_ ( .D(
        mem_stage_inst_dmem_n3145), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__5_ ( .D(
        mem_stage_inst_dmem_n3146), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__6_ ( .D(
        mem_stage_inst_dmem_n3147), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__7_ ( .D(
        mem_stage_inst_dmem_n3148), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__8_ ( .D(
        mem_stage_inst_dmem_n3149), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__9_ ( .D(
        mem_stage_inst_dmem_n3150), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__10_ ( .D(
        mem_stage_inst_dmem_n3151), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__11_ ( .D(
        mem_stage_inst_dmem_n3152), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__12_ ( .D(
        mem_stage_inst_dmem_n3153), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__13_ ( .D(
        mem_stage_inst_dmem_n3154), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__14_ ( .D(
        mem_stage_inst_dmem_n3155), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_161__15_ ( .D(
        mem_stage_inst_dmem_n3156), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_161__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__0_ ( .D(
        mem_stage_inst_dmem_n3205), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__1_ ( .D(
        mem_stage_inst_dmem_n3206), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__2_ ( .D(
        mem_stage_inst_dmem_n3207), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__3_ ( .D(
        mem_stage_inst_dmem_n3208), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__4_ ( .D(
        mem_stage_inst_dmem_n3209), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__5_ ( .D(
        mem_stage_inst_dmem_n3210), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__6_ ( .D(
        mem_stage_inst_dmem_n3211), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__7_ ( .D(
        mem_stage_inst_dmem_n3212), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__8_ ( .D(
        mem_stage_inst_dmem_n3213), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__9_ ( .D(
        mem_stage_inst_dmem_n3214), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__10_ ( .D(
        mem_stage_inst_dmem_n3215), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__11_ ( .D(
        mem_stage_inst_dmem_n3216), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__12_ ( .D(
        mem_stage_inst_dmem_n3217), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__13_ ( .D(
        mem_stage_inst_dmem_n3218), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__14_ ( .D(
        mem_stage_inst_dmem_n3219), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_165__15_ ( .D(
        mem_stage_inst_dmem_n3220), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_165__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__0_ ( .D(
        mem_stage_inst_dmem_n3269), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__1_ ( .D(
        mem_stage_inst_dmem_n3270), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__2_ ( .D(
        mem_stage_inst_dmem_n3271), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__3_ ( .D(
        mem_stage_inst_dmem_n3272), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__4_ ( .D(
        mem_stage_inst_dmem_n3273), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__5_ ( .D(
        mem_stage_inst_dmem_n3274), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__6_ ( .D(
        mem_stage_inst_dmem_n3275), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__7_ ( .D(
        mem_stage_inst_dmem_n3276), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__8_ ( .D(
        mem_stage_inst_dmem_n3277), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__9_ ( .D(
        mem_stage_inst_dmem_n3278), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__10_ ( .D(
        mem_stage_inst_dmem_n3279), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__11_ ( .D(
        mem_stage_inst_dmem_n3280), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__12_ ( .D(
        mem_stage_inst_dmem_n3281), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__13_ ( .D(
        mem_stage_inst_dmem_n3282), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__14_ ( .D(
        mem_stage_inst_dmem_n3283), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_169__15_ ( .D(
        mem_stage_inst_dmem_n3284), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_169__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__0_ ( .D(
        mem_stage_inst_dmem_n3333), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__1_ ( .D(
        mem_stage_inst_dmem_n3334), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__2_ ( .D(
        mem_stage_inst_dmem_n3335), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__3_ ( .D(
        mem_stage_inst_dmem_n3336), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__4_ ( .D(
        mem_stage_inst_dmem_n3337), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__5_ ( .D(
        mem_stage_inst_dmem_n3338), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__6_ ( .D(
        mem_stage_inst_dmem_n3339), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__7_ ( .D(
        mem_stage_inst_dmem_n3340), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__8_ ( .D(
        mem_stage_inst_dmem_n3341), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__9_ ( .D(
        mem_stage_inst_dmem_n3342), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__10_ ( .D(
        mem_stage_inst_dmem_n3343), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__11_ ( .D(
        mem_stage_inst_dmem_n3344), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__12_ ( .D(
        mem_stage_inst_dmem_n3345), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__13_ ( .D(
        mem_stage_inst_dmem_n3346), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__14_ ( .D(
        mem_stage_inst_dmem_n3347), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_173__15_ ( .D(
        mem_stage_inst_dmem_n3348), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_173__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__0_ ( .D(
        mem_stage_inst_dmem_n3397), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__1_ ( .D(
        mem_stage_inst_dmem_n3398), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__2_ ( .D(
        mem_stage_inst_dmem_n3399), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__3_ ( .D(
        mem_stage_inst_dmem_n3400), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__4_ ( .D(
        mem_stage_inst_dmem_n3401), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__5_ ( .D(
        mem_stage_inst_dmem_n3402), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__6_ ( .D(
        mem_stage_inst_dmem_n3403), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__7_ ( .D(
        mem_stage_inst_dmem_n3404), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__8_ ( .D(
        mem_stage_inst_dmem_n3405), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__9_ ( .D(
        mem_stage_inst_dmem_n3406), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__10_ ( .D(
        mem_stage_inst_dmem_n3407), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__11_ ( .D(
        mem_stage_inst_dmem_n3408), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__12_ ( .D(
        mem_stage_inst_dmem_n3409), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__13_ ( .D(
        mem_stage_inst_dmem_n3410), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__14_ ( .D(
        mem_stage_inst_dmem_n3411), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_177__15_ ( .D(
        mem_stage_inst_dmem_n3412), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_177__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__0_ ( .D(
        mem_stage_inst_dmem_n3461), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__1_ ( .D(
        mem_stage_inst_dmem_n3462), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__2_ ( .D(
        mem_stage_inst_dmem_n3463), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__3_ ( .D(
        mem_stage_inst_dmem_n3464), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__4_ ( .D(
        mem_stage_inst_dmem_n3465), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__5_ ( .D(
        mem_stage_inst_dmem_n3466), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__6_ ( .D(
        mem_stage_inst_dmem_n3467), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__7_ ( .D(
        mem_stage_inst_dmem_n3468), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__8_ ( .D(
        mem_stage_inst_dmem_n3469), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__9_ ( .D(
        mem_stage_inst_dmem_n3470), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__10_ ( .D(
        mem_stage_inst_dmem_n3471), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__11_ ( .D(
        mem_stage_inst_dmem_n3472), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__12_ ( .D(
        mem_stage_inst_dmem_n3473), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__13_ ( .D(
        mem_stage_inst_dmem_n3474), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__14_ ( .D(
        mem_stage_inst_dmem_n3475), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_181__15_ ( .D(
        mem_stage_inst_dmem_n3476), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_181__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__0_ ( .D(
        mem_stage_inst_dmem_n3525), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__1_ ( .D(
        mem_stage_inst_dmem_n3526), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__2_ ( .D(
        mem_stage_inst_dmem_n3527), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__3_ ( .D(
        mem_stage_inst_dmem_n3528), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__4_ ( .D(
        mem_stage_inst_dmem_n3529), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__5_ ( .D(
        mem_stage_inst_dmem_n3530), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__6_ ( .D(
        mem_stage_inst_dmem_n3531), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__7_ ( .D(
        mem_stage_inst_dmem_n3532), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__8_ ( .D(
        mem_stage_inst_dmem_n3533), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__9_ ( .D(
        mem_stage_inst_dmem_n3534), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__10_ ( .D(
        mem_stage_inst_dmem_n3535), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__11_ ( .D(
        mem_stage_inst_dmem_n3536), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__12_ ( .D(
        mem_stage_inst_dmem_n3537), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__13_ ( .D(
        mem_stage_inst_dmem_n3538), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__14_ ( .D(
        mem_stage_inst_dmem_n3539), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_185__15_ ( .D(
        mem_stage_inst_dmem_n3540), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_185__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__0_ ( .D(
        mem_stage_inst_dmem_n3589), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__1_ ( .D(
        mem_stage_inst_dmem_n3590), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__2_ ( .D(
        mem_stage_inst_dmem_n3591), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__3_ ( .D(
        mem_stage_inst_dmem_n3592), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__4_ ( .D(
        mem_stage_inst_dmem_n3593), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__5_ ( .D(
        mem_stage_inst_dmem_n3594), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__6_ ( .D(
        mem_stage_inst_dmem_n3595), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__7_ ( .D(
        mem_stage_inst_dmem_n3596), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__8_ ( .D(
        mem_stage_inst_dmem_n3597), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__9_ ( .D(
        mem_stage_inst_dmem_n3598), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__10_ ( .D(
        mem_stage_inst_dmem_n3599), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__11_ ( .D(
        mem_stage_inst_dmem_n3600), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__12_ ( .D(
        mem_stage_inst_dmem_n3601), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__13_ ( .D(
        mem_stage_inst_dmem_n3602), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__14_ ( .D(
        mem_stage_inst_dmem_n3603), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_189__15_ ( .D(
        mem_stage_inst_dmem_n3604), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_189__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__0_ ( .D(
        mem_stage_inst_dmem_n3653), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__1_ ( .D(
        mem_stage_inst_dmem_n3654), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__2_ ( .D(
        mem_stage_inst_dmem_n3655), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__3_ ( .D(
        mem_stage_inst_dmem_n3656), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__4_ ( .D(
        mem_stage_inst_dmem_n3657), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__5_ ( .D(
        mem_stage_inst_dmem_n3658), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__6_ ( .D(
        mem_stage_inst_dmem_n3659), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__7_ ( .D(
        mem_stage_inst_dmem_n3660), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__8_ ( .D(
        mem_stage_inst_dmem_n3661), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__9_ ( .D(
        mem_stage_inst_dmem_n3662), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__10_ ( .D(
        mem_stage_inst_dmem_n3663), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__11_ ( .D(
        mem_stage_inst_dmem_n3664), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__12_ ( .D(
        mem_stage_inst_dmem_n3665), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__13_ ( .D(
        mem_stage_inst_dmem_n3666), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__14_ ( .D(
        mem_stage_inst_dmem_n3667), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_193__15_ ( .D(
        mem_stage_inst_dmem_n3668), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_193__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__0_ ( .D(
        mem_stage_inst_dmem_n3717), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__1_ ( .D(
        mem_stage_inst_dmem_n3718), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__2_ ( .D(
        mem_stage_inst_dmem_n3719), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__3_ ( .D(
        mem_stage_inst_dmem_n3720), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__4_ ( .D(
        mem_stage_inst_dmem_n3721), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__5_ ( .D(
        mem_stage_inst_dmem_n3722), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__6_ ( .D(
        mem_stage_inst_dmem_n3723), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__7_ ( .D(
        mem_stage_inst_dmem_n3724), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__8_ ( .D(
        mem_stage_inst_dmem_n3725), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__9_ ( .D(
        mem_stage_inst_dmem_n3726), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__10_ ( .D(
        mem_stage_inst_dmem_n3727), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__11_ ( .D(
        mem_stage_inst_dmem_n3728), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__12_ ( .D(
        mem_stage_inst_dmem_n3729), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__13_ ( .D(
        mem_stage_inst_dmem_n3730), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__14_ ( .D(
        mem_stage_inst_dmem_n3731), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_197__15_ ( .D(
        mem_stage_inst_dmem_n3732), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_197__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__0_ ( .D(
        mem_stage_inst_dmem_n3781), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__1_ ( .D(
        mem_stage_inst_dmem_n3782), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__2_ ( .D(
        mem_stage_inst_dmem_n3783), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__3_ ( .D(
        mem_stage_inst_dmem_n3784), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__4_ ( .D(
        mem_stage_inst_dmem_n3785), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__5_ ( .D(
        mem_stage_inst_dmem_n3786), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__6_ ( .D(
        mem_stage_inst_dmem_n3787), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__7_ ( .D(
        mem_stage_inst_dmem_n3788), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__8_ ( .D(
        mem_stage_inst_dmem_n3789), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__9_ ( .D(
        mem_stage_inst_dmem_n3790), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__10_ ( .D(
        mem_stage_inst_dmem_n3791), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__11_ ( .D(
        mem_stage_inst_dmem_n3792), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__12_ ( .D(
        mem_stage_inst_dmem_n3793), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__13_ ( .D(
        mem_stage_inst_dmem_n3794), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__14_ ( .D(
        mem_stage_inst_dmem_n3795), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_201__15_ ( .D(
        mem_stage_inst_dmem_n3796), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_201__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__0_ ( .D(
        mem_stage_inst_dmem_n3845), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__1_ ( .D(
        mem_stage_inst_dmem_n3846), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__2_ ( .D(
        mem_stage_inst_dmem_n3847), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__3_ ( .D(
        mem_stage_inst_dmem_n3848), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__4_ ( .D(
        mem_stage_inst_dmem_n3849), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__5_ ( .D(
        mem_stage_inst_dmem_n3850), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__6_ ( .D(
        mem_stage_inst_dmem_n3851), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__7_ ( .D(
        mem_stage_inst_dmem_n3852), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__8_ ( .D(
        mem_stage_inst_dmem_n3853), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__9_ ( .D(
        mem_stage_inst_dmem_n3854), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__10_ ( .D(
        mem_stage_inst_dmem_n3855), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__11_ ( .D(
        mem_stage_inst_dmem_n3856), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__12_ ( .D(
        mem_stage_inst_dmem_n3857), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__13_ ( .D(
        mem_stage_inst_dmem_n3858), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__14_ ( .D(
        mem_stage_inst_dmem_n3859), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_205__15_ ( .D(
        mem_stage_inst_dmem_n3860), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_205__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__0_ ( .D(
        mem_stage_inst_dmem_n3909), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__1_ ( .D(
        mem_stage_inst_dmem_n3910), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__2_ ( .D(
        mem_stage_inst_dmem_n3911), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__3_ ( .D(
        mem_stage_inst_dmem_n3912), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__4_ ( .D(
        mem_stage_inst_dmem_n3913), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__5_ ( .D(
        mem_stage_inst_dmem_n3914), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__6_ ( .D(
        mem_stage_inst_dmem_n3915), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__7_ ( .D(
        mem_stage_inst_dmem_n3916), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__8_ ( .D(
        mem_stage_inst_dmem_n3917), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__9_ ( .D(
        mem_stage_inst_dmem_n3918), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__10_ ( .D(
        mem_stage_inst_dmem_n3919), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__11_ ( .D(
        mem_stage_inst_dmem_n3920), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__12_ ( .D(
        mem_stage_inst_dmem_n3921), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__13_ ( .D(
        mem_stage_inst_dmem_n3922), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__14_ ( .D(
        mem_stage_inst_dmem_n3923), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_209__15_ ( .D(
        mem_stage_inst_dmem_n3924), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_209__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__0_ ( .D(
        mem_stage_inst_dmem_n3973), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__1_ ( .D(
        mem_stage_inst_dmem_n3974), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__2_ ( .D(
        mem_stage_inst_dmem_n3975), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__3_ ( .D(
        mem_stage_inst_dmem_n3976), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__4_ ( .D(
        mem_stage_inst_dmem_n3977), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__5_ ( .D(
        mem_stage_inst_dmem_n3978), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__6_ ( .D(
        mem_stage_inst_dmem_n3979), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__7_ ( .D(
        mem_stage_inst_dmem_n3980), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__8_ ( .D(
        mem_stage_inst_dmem_n3981), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__9_ ( .D(
        mem_stage_inst_dmem_n3982), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__10_ ( .D(
        mem_stage_inst_dmem_n3983), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__11_ ( .D(
        mem_stage_inst_dmem_n3984), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__12_ ( .D(
        mem_stage_inst_dmem_n3985), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__13_ ( .D(
        mem_stage_inst_dmem_n3986), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__14_ ( .D(
        mem_stage_inst_dmem_n3987), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_213__15_ ( .D(
        mem_stage_inst_dmem_n3988), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_213__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__0_ ( .D(
        mem_stage_inst_dmem_n4037), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__1_ ( .D(
        mem_stage_inst_dmem_n4038), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__2_ ( .D(
        mem_stage_inst_dmem_n4039), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__3_ ( .D(
        mem_stage_inst_dmem_n4040), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__4_ ( .D(
        mem_stage_inst_dmem_n4041), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__5_ ( .D(
        mem_stage_inst_dmem_n4042), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__6_ ( .D(
        mem_stage_inst_dmem_n4043), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__7_ ( .D(
        mem_stage_inst_dmem_n4044), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__8_ ( .D(
        mem_stage_inst_dmem_n4045), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__9_ ( .D(
        mem_stage_inst_dmem_n4046), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__10_ ( .D(
        mem_stage_inst_dmem_n4047), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__11_ ( .D(
        mem_stage_inst_dmem_n4048), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__12_ ( .D(
        mem_stage_inst_dmem_n4049), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__13_ ( .D(
        mem_stage_inst_dmem_n4050), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__14_ ( .D(
        mem_stage_inst_dmem_n4051), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_217__15_ ( .D(
        mem_stage_inst_dmem_n4052), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_217__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__0_ ( .D(
        mem_stage_inst_dmem_n4101), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__1_ ( .D(
        mem_stage_inst_dmem_n4102), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__2_ ( .D(
        mem_stage_inst_dmem_n4103), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__3_ ( .D(
        mem_stage_inst_dmem_n4104), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__4_ ( .D(
        mem_stage_inst_dmem_n4105), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__5_ ( .D(
        mem_stage_inst_dmem_n4106), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__6_ ( .D(
        mem_stage_inst_dmem_n4107), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__7_ ( .D(
        mem_stage_inst_dmem_n4108), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__8_ ( .D(
        mem_stage_inst_dmem_n4109), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__9_ ( .D(
        mem_stage_inst_dmem_n4110), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__10_ ( .D(
        mem_stage_inst_dmem_n4111), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__11_ ( .D(
        mem_stage_inst_dmem_n4112), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__12_ ( .D(
        mem_stage_inst_dmem_n4113), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__13_ ( .D(
        mem_stage_inst_dmem_n4114), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__14_ ( .D(
        mem_stage_inst_dmem_n4115), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_221__15_ ( .D(
        mem_stage_inst_dmem_n4116), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_221__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__0_ ( .D(
        mem_stage_inst_dmem_n4165), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__1_ ( .D(
        mem_stage_inst_dmem_n4166), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__2_ ( .D(
        mem_stage_inst_dmem_n4167), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__3_ ( .D(
        mem_stage_inst_dmem_n4168), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__4_ ( .D(
        mem_stage_inst_dmem_n4169), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__5_ ( .D(
        mem_stage_inst_dmem_n4170), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__6_ ( .D(
        mem_stage_inst_dmem_n4171), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__7_ ( .D(
        mem_stage_inst_dmem_n4172), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__8_ ( .D(
        mem_stage_inst_dmem_n4173), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__9_ ( .D(
        mem_stage_inst_dmem_n4174), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__10_ ( .D(
        mem_stage_inst_dmem_n4175), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__11_ ( .D(
        mem_stage_inst_dmem_n4176), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__12_ ( .D(
        mem_stage_inst_dmem_n4177), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__13_ ( .D(
        mem_stage_inst_dmem_n4178), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__14_ ( .D(
        mem_stage_inst_dmem_n4179), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_225__15_ ( .D(
        mem_stage_inst_dmem_n4180), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_225__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__0_ ( .D(
        mem_stage_inst_dmem_n4229), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__1_ ( .D(
        mem_stage_inst_dmem_n4230), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__2_ ( .D(
        mem_stage_inst_dmem_n4231), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__3_ ( .D(
        mem_stage_inst_dmem_n4232), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__4_ ( .D(
        mem_stage_inst_dmem_n4233), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__5_ ( .D(
        mem_stage_inst_dmem_n4234), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__6_ ( .D(
        mem_stage_inst_dmem_n4235), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__7_ ( .D(
        mem_stage_inst_dmem_n4236), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__8_ ( .D(
        mem_stage_inst_dmem_n4237), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__9_ ( .D(
        mem_stage_inst_dmem_n4238), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__10_ ( .D(
        mem_stage_inst_dmem_n4239), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__11_ ( .D(
        mem_stage_inst_dmem_n4240), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__12_ ( .D(
        mem_stage_inst_dmem_n4241), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__13_ ( .D(
        mem_stage_inst_dmem_n4242), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__14_ ( .D(
        mem_stage_inst_dmem_n4243), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_229__15_ ( .D(
        mem_stage_inst_dmem_n4244), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_229__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__0_ ( .D(
        mem_stage_inst_dmem_n4293), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__1_ ( .D(
        mem_stage_inst_dmem_n4294), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__2_ ( .D(
        mem_stage_inst_dmem_n4295), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__3_ ( .D(
        mem_stage_inst_dmem_n4296), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__4_ ( .D(
        mem_stage_inst_dmem_n4297), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__5_ ( .D(
        mem_stage_inst_dmem_n4298), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__6_ ( .D(
        mem_stage_inst_dmem_n4299), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__7_ ( .D(
        mem_stage_inst_dmem_n4300), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__8_ ( .D(
        mem_stage_inst_dmem_n4301), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__9_ ( .D(
        mem_stage_inst_dmem_n4302), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__10_ ( .D(
        mem_stage_inst_dmem_n4303), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__11_ ( .D(
        mem_stage_inst_dmem_n4304), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__12_ ( .D(
        mem_stage_inst_dmem_n4305), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__13_ ( .D(
        mem_stage_inst_dmem_n4306), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__14_ ( .D(
        mem_stage_inst_dmem_n4307), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_233__15_ ( .D(
        mem_stage_inst_dmem_n4308), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_233__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__0_ ( .D(
        mem_stage_inst_dmem_n4357), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__1_ ( .D(
        mem_stage_inst_dmem_n4358), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__2_ ( .D(
        mem_stage_inst_dmem_n4359), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__3_ ( .D(
        mem_stage_inst_dmem_n4360), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__4_ ( .D(
        mem_stage_inst_dmem_n4361), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__5_ ( .D(
        mem_stage_inst_dmem_n4362), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__6_ ( .D(
        mem_stage_inst_dmem_n4363), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__7_ ( .D(
        mem_stage_inst_dmem_n4364), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__8_ ( .D(
        mem_stage_inst_dmem_n4365), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__9_ ( .D(
        mem_stage_inst_dmem_n4366), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__10_ ( .D(
        mem_stage_inst_dmem_n4367), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__11_ ( .D(
        mem_stage_inst_dmem_n4368), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__12_ ( .D(
        mem_stage_inst_dmem_n4369), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__13_ ( .D(
        mem_stage_inst_dmem_n4370), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__14_ ( .D(
        mem_stage_inst_dmem_n4371), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_237__15_ ( .D(
        mem_stage_inst_dmem_n4372), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_237__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__0_ ( .D(
        mem_stage_inst_dmem_n4421), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__1_ ( .D(
        mem_stage_inst_dmem_n4422), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__2_ ( .D(
        mem_stage_inst_dmem_n4423), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__3_ ( .D(
        mem_stage_inst_dmem_n4424), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__4_ ( .D(
        mem_stage_inst_dmem_n4425), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__5_ ( .D(
        mem_stage_inst_dmem_n4426), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__6_ ( .D(
        mem_stage_inst_dmem_n4427), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__7_ ( .D(
        mem_stage_inst_dmem_n4428), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__8_ ( .D(
        mem_stage_inst_dmem_n4429), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__9_ ( .D(
        mem_stage_inst_dmem_n4430), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__10_ ( .D(
        mem_stage_inst_dmem_n4431), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__11_ ( .D(
        mem_stage_inst_dmem_n4432), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__12_ ( .D(
        mem_stage_inst_dmem_n4433), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__13_ ( .D(
        mem_stage_inst_dmem_n4434), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__14_ ( .D(
        mem_stage_inst_dmem_n4435), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_241__15_ ( .D(
        mem_stage_inst_dmem_n4436), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_241__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__0_ ( .D(
        mem_stage_inst_dmem_n4485), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__1_ ( .D(
        mem_stage_inst_dmem_n4486), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__2_ ( .D(
        mem_stage_inst_dmem_n4487), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__3_ ( .D(
        mem_stage_inst_dmem_n4488), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__4_ ( .D(
        mem_stage_inst_dmem_n4489), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__5_ ( .D(
        mem_stage_inst_dmem_n4490), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__6_ ( .D(
        mem_stage_inst_dmem_n4491), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__7_ ( .D(
        mem_stage_inst_dmem_n4492), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__8_ ( .D(
        mem_stage_inst_dmem_n4493), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__9_ ( .D(
        mem_stage_inst_dmem_n4494), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__10_ ( .D(
        mem_stage_inst_dmem_n4495), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__11_ ( .D(
        mem_stage_inst_dmem_n4496), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__12_ ( .D(
        mem_stage_inst_dmem_n4497), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__13_ ( .D(
        mem_stage_inst_dmem_n4498), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__14_ ( .D(
        mem_stage_inst_dmem_n4499), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_245__15_ ( .D(
        mem_stage_inst_dmem_n4500), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_245__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__0_ ( .D(
        mem_stage_inst_dmem_n4549), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__1_ ( .D(
        mem_stage_inst_dmem_n4550), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__2_ ( .D(
        mem_stage_inst_dmem_n4551), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__3_ ( .D(
        mem_stage_inst_dmem_n4552), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__4_ ( .D(
        mem_stage_inst_dmem_n4553), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__5_ ( .D(
        mem_stage_inst_dmem_n4554), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__6_ ( .D(
        mem_stage_inst_dmem_n4555), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__7_ ( .D(
        mem_stage_inst_dmem_n4556), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__8_ ( .D(
        mem_stage_inst_dmem_n4557), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__9_ ( .D(
        mem_stage_inst_dmem_n4558), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__10_ ( .D(
        mem_stage_inst_dmem_n4559), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__11_ ( .D(
        mem_stage_inst_dmem_n4560), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__12_ ( .D(
        mem_stage_inst_dmem_n4561), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__13_ ( .D(
        mem_stage_inst_dmem_n4562), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__14_ ( .D(
        mem_stage_inst_dmem_n4563), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_249__15_ ( .D(
        mem_stage_inst_dmem_n4564), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_249__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__0_ ( .D(
        mem_stage_inst_dmem_n4613), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__1_ ( .D(
        mem_stage_inst_dmem_n4614), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__2_ ( .D(
        mem_stage_inst_dmem_n4615), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__3_ ( .D(
        mem_stage_inst_dmem_n4616), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__4_ ( .D(
        mem_stage_inst_dmem_n4617), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__5_ ( .D(
        mem_stage_inst_dmem_n4618), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__6_ ( .D(
        mem_stage_inst_dmem_n4619), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__7_ ( .D(
        mem_stage_inst_dmem_n4620), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__8_ ( .D(
        mem_stage_inst_dmem_n4621), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__9_ ( .D(
        mem_stage_inst_dmem_n4622), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__10_ ( .D(
        mem_stage_inst_dmem_n4623), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__11_ ( .D(
        mem_stage_inst_dmem_n4624), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__12_ ( .D(
        mem_stage_inst_dmem_n4625), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__13_ ( .D(
        mem_stage_inst_dmem_n4626), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__14_ ( .D(
        mem_stage_inst_dmem_n4627), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_253__15_ ( .D(
        mem_stage_inst_dmem_n4628), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_253__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__0_ ( .D(
        mem_stage_inst_dmem_n613), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__1_ ( .D(
        mem_stage_inst_dmem_n614), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__2_ ( .D(
        mem_stage_inst_dmem_n615), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__3_ ( .D(
        mem_stage_inst_dmem_n616), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__4_ ( .D(
        mem_stage_inst_dmem_n617), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__5_ ( .D(
        mem_stage_inst_dmem_n618), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__6_ ( .D(
        mem_stage_inst_dmem_n619), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__7_ ( .D(
        mem_stage_inst_dmem_n620), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__8_ ( .D(
        mem_stage_inst_dmem_n621), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__9_ ( .D(
        mem_stage_inst_dmem_n622), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__10_ ( .D(
        mem_stage_inst_dmem_n623), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__11_ ( .D(
        mem_stage_inst_dmem_n624), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__12_ ( .D(
        mem_stage_inst_dmem_n625), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__13_ ( .D(
        mem_stage_inst_dmem_n626), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__14_ ( .D(
        mem_stage_inst_dmem_n627), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_3__15_ ( .D(
        mem_stage_inst_dmem_n628), .CK(clk), .Q(mem_stage_inst_dmem_ram_3__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__0_ ( .D(
        mem_stage_inst_dmem_n677), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__0_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__1_ ( .D(
        mem_stage_inst_dmem_n678), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__1_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__2_ ( .D(
        mem_stage_inst_dmem_n679), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__2_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__3_ ( .D(
        mem_stage_inst_dmem_n680), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__3_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__4_ ( .D(
        mem_stage_inst_dmem_n681), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__4_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__5_ ( .D(
        mem_stage_inst_dmem_n682), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__5_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__6_ ( .D(
        mem_stage_inst_dmem_n683), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__6_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__7_ ( .D(
        mem_stage_inst_dmem_n684), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__7_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__8_ ( .D(
        mem_stage_inst_dmem_n685), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__8_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__9_ ( .D(
        mem_stage_inst_dmem_n686), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__9_)
         );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__10_ ( .D(
        mem_stage_inst_dmem_n687), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__11_ ( .D(
        mem_stage_inst_dmem_n688), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__12_ ( .D(
        mem_stage_inst_dmem_n689), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__13_ ( .D(
        mem_stage_inst_dmem_n690), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__14_ ( .D(
        mem_stage_inst_dmem_n691), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_7__15_ ( .D(
        mem_stage_inst_dmem_n692), .CK(clk), .Q(mem_stage_inst_dmem_ram_7__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__0_ ( .D(
        mem_stage_inst_dmem_n741), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__1_ ( .D(
        mem_stage_inst_dmem_n742), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__2_ ( .D(
        mem_stage_inst_dmem_n743), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__3_ ( .D(
        mem_stage_inst_dmem_n744), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__4_ ( .D(
        mem_stage_inst_dmem_n745), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__5_ ( .D(
        mem_stage_inst_dmem_n746), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__6_ ( .D(
        mem_stage_inst_dmem_n747), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__7_ ( .D(
        mem_stage_inst_dmem_n748), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__8_ ( .D(
        mem_stage_inst_dmem_n749), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__9_ ( .D(
        mem_stage_inst_dmem_n750), .CK(clk), .Q(mem_stage_inst_dmem_ram_11__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__10_ ( .D(
        mem_stage_inst_dmem_n751), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_11__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__11_ ( .D(
        mem_stage_inst_dmem_n752), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_11__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__12_ ( .D(
        mem_stage_inst_dmem_n753), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_11__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__13_ ( .D(
        mem_stage_inst_dmem_n754), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_11__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__14_ ( .D(
        mem_stage_inst_dmem_n755), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_11__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_11__15_ ( .D(
        mem_stage_inst_dmem_n756), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_11__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__0_ ( .D(
        mem_stage_inst_dmem_n805), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__1_ ( .D(
        mem_stage_inst_dmem_n806), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__2_ ( .D(
        mem_stage_inst_dmem_n807), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__3_ ( .D(
        mem_stage_inst_dmem_n808), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__4_ ( .D(
        mem_stage_inst_dmem_n809), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__5_ ( .D(
        mem_stage_inst_dmem_n810), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__6_ ( .D(
        mem_stage_inst_dmem_n811), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__7_ ( .D(
        mem_stage_inst_dmem_n812), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__8_ ( .D(
        mem_stage_inst_dmem_n813), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__9_ ( .D(
        mem_stage_inst_dmem_n814), .CK(clk), .Q(mem_stage_inst_dmem_ram_15__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__10_ ( .D(
        mem_stage_inst_dmem_n815), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_15__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__11_ ( .D(
        mem_stage_inst_dmem_n816), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_15__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__12_ ( .D(
        mem_stage_inst_dmem_n817), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_15__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__13_ ( .D(
        mem_stage_inst_dmem_n818), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_15__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__14_ ( .D(
        mem_stage_inst_dmem_n819), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_15__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_15__15_ ( .D(
        mem_stage_inst_dmem_n820), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_15__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__0_ ( .D(
        mem_stage_inst_dmem_n869), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__1_ ( .D(
        mem_stage_inst_dmem_n870), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__2_ ( .D(
        mem_stage_inst_dmem_n871), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__3_ ( .D(
        mem_stage_inst_dmem_n872), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__4_ ( .D(
        mem_stage_inst_dmem_n873), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__5_ ( .D(
        mem_stage_inst_dmem_n874), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__6_ ( .D(
        mem_stage_inst_dmem_n875), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__7_ ( .D(
        mem_stage_inst_dmem_n876), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__8_ ( .D(
        mem_stage_inst_dmem_n877), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__9_ ( .D(
        mem_stage_inst_dmem_n878), .CK(clk), .Q(mem_stage_inst_dmem_ram_19__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__10_ ( .D(
        mem_stage_inst_dmem_n879), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_19__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__11_ ( .D(
        mem_stage_inst_dmem_n880), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_19__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__12_ ( .D(
        mem_stage_inst_dmem_n881), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_19__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__13_ ( .D(
        mem_stage_inst_dmem_n882), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_19__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__14_ ( .D(
        mem_stage_inst_dmem_n883), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_19__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_19__15_ ( .D(
        mem_stage_inst_dmem_n884), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_19__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__0_ ( .D(
        mem_stage_inst_dmem_n933), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__1_ ( .D(
        mem_stage_inst_dmem_n934), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__2_ ( .D(
        mem_stage_inst_dmem_n935), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__3_ ( .D(
        mem_stage_inst_dmem_n936), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__4_ ( .D(
        mem_stage_inst_dmem_n937), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__5_ ( .D(
        mem_stage_inst_dmem_n938), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__6_ ( .D(
        mem_stage_inst_dmem_n939), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__7_ ( .D(
        mem_stage_inst_dmem_n940), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__8_ ( .D(
        mem_stage_inst_dmem_n941), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__9_ ( .D(
        mem_stage_inst_dmem_n942), .CK(clk), .Q(mem_stage_inst_dmem_ram_23__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__10_ ( .D(
        mem_stage_inst_dmem_n943), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_23__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__11_ ( .D(
        mem_stage_inst_dmem_n944), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_23__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__12_ ( .D(
        mem_stage_inst_dmem_n945), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_23__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__13_ ( .D(
        mem_stage_inst_dmem_n946), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_23__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__14_ ( .D(
        mem_stage_inst_dmem_n947), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_23__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_23__15_ ( .D(
        mem_stage_inst_dmem_n948), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_23__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__0_ ( .D(
        mem_stage_inst_dmem_n997), .CK(clk), .Q(mem_stage_inst_dmem_ram_27__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__1_ ( .D(
        mem_stage_inst_dmem_n998), .CK(clk), .Q(mem_stage_inst_dmem_ram_27__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__2_ ( .D(
        mem_stage_inst_dmem_n999), .CK(clk), .Q(mem_stage_inst_dmem_ram_27__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__3_ ( .D(
        mem_stage_inst_dmem_n1000), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__4_ ( .D(
        mem_stage_inst_dmem_n1001), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__5_ ( .D(
        mem_stage_inst_dmem_n1002), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__6_ ( .D(
        mem_stage_inst_dmem_n1003), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__7_ ( .D(
        mem_stage_inst_dmem_n1004), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__8_ ( .D(
        mem_stage_inst_dmem_n1005), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__9_ ( .D(
        mem_stage_inst_dmem_n1006), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__10_ ( .D(
        mem_stage_inst_dmem_n1007), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__11_ ( .D(
        mem_stage_inst_dmem_n1008), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__12_ ( .D(
        mem_stage_inst_dmem_n1009), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__13_ ( .D(
        mem_stage_inst_dmem_n1010), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__14_ ( .D(
        mem_stage_inst_dmem_n1011), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_27__15_ ( .D(
        mem_stage_inst_dmem_n1012), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_27__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__0_ ( .D(
        mem_stage_inst_dmem_n1061), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__1_ ( .D(
        mem_stage_inst_dmem_n1062), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__2_ ( .D(
        mem_stage_inst_dmem_n1063), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__3_ ( .D(
        mem_stage_inst_dmem_n1064), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__4_ ( .D(
        mem_stage_inst_dmem_n1065), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__5_ ( .D(
        mem_stage_inst_dmem_n1066), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__6_ ( .D(
        mem_stage_inst_dmem_n1067), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__7_ ( .D(
        mem_stage_inst_dmem_n1068), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__8_ ( .D(
        mem_stage_inst_dmem_n1069), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__9_ ( .D(
        mem_stage_inst_dmem_n1070), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__10_ ( .D(
        mem_stage_inst_dmem_n1071), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__11_ ( .D(
        mem_stage_inst_dmem_n1072), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__12_ ( .D(
        mem_stage_inst_dmem_n1073), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__13_ ( .D(
        mem_stage_inst_dmem_n1074), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__14_ ( .D(
        mem_stage_inst_dmem_n1075), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_31__15_ ( .D(
        mem_stage_inst_dmem_n1076), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_31__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__0_ ( .D(
        mem_stage_inst_dmem_n1125), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__1_ ( .D(
        mem_stage_inst_dmem_n1126), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__2_ ( .D(
        mem_stage_inst_dmem_n1127), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__3_ ( .D(
        mem_stage_inst_dmem_n1128), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__4_ ( .D(
        mem_stage_inst_dmem_n1129), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__5_ ( .D(
        mem_stage_inst_dmem_n1130), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__6_ ( .D(
        mem_stage_inst_dmem_n1131), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__7_ ( .D(
        mem_stage_inst_dmem_n1132), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__8_ ( .D(
        mem_stage_inst_dmem_n1133), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__9_ ( .D(
        mem_stage_inst_dmem_n1134), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__10_ ( .D(
        mem_stage_inst_dmem_n1135), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__11_ ( .D(
        mem_stage_inst_dmem_n1136), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__12_ ( .D(
        mem_stage_inst_dmem_n1137), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__13_ ( .D(
        mem_stage_inst_dmem_n1138), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__14_ ( .D(
        mem_stage_inst_dmem_n1139), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_35__15_ ( .D(
        mem_stage_inst_dmem_n1140), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_35__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__0_ ( .D(
        mem_stage_inst_dmem_n1189), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__1_ ( .D(
        mem_stage_inst_dmem_n1190), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__2_ ( .D(
        mem_stage_inst_dmem_n1191), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__3_ ( .D(
        mem_stage_inst_dmem_n1192), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__4_ ( .D(
        mem_stage_inst_dmem_n1193), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__5_ ( .D(
        mem_stage_inst_dmem_n1194), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__6_ ( .D(
        mem_stage_inst_dmem_n1195), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__7_ ( .D(
        mem_stage_inst_dmem_n1196), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__8_ ( .D(
        mem_stage_inst_dmem_n1197), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__9_ ( .D(
        mem_stage_inst_dmem_n1198), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__10_ ( .D(
        mem_stage_inst_dmem_n1199), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__11_ ( .D(
        mem_stage_inst_dmem_n1200), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__12_ ( .D(
        mem_stage_inst_dmem_n1201), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__13_ ( .D(
        mem_stage_inst_dmem_n1202), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__14_ ( .D(
        mem_stage_inst_dmem_n1203), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_39__15_ ( .D(
        mem_stage_inst_dmem_n1204), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_39__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__0_ ( .D(
        mem_stage_inst_dmem_n1253), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__1_ ( .D(
        mem_stage_inst_dmem_n1254), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__2_ ( .D(
        mem_stage_inst_dmem_n1255), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__3_ ( .D(
        mem_stage_inst_dmem_n1256), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__4_ ( .D(
        mem_stage_inst_dmem_n1257), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__5_ ( .D(
        mem_stage_inst_dmem_n1258), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__6_ ( .D(
        mem_stage_inst_dmem_n1259), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__7_ ( .D(
        mem_stage_inst_dmem_n1260), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__8_ ( .D(
        mem_stage_inst_dmem_n1261), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__9_ ( .D(
        mem_stage_inst_dmem_n1262), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__10_ ( .D(
        mem_stage_inst_dmem_n1263), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__11_ ( .D(
        mem_stage_inst_dmem_n1264), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__12_ ( .D(
        mem_stage_inst_dmem_n1265), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__13_ ( .D(
        mem_stage_inst_dmem_n1266), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__14_ ( .D(
        mem_stage_inst_dmem_n1267), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_43__15_ ( .D(
        mem_stage_inst_dmem_n1268), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_43__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__0_ ( .D(
        mem_stage_inst_dmem_n1317), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__1_ ( .D(
        mem_stage_inst_dmem_n1318), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__2_ ( .D(
        mem_stage_inst_dmem_n1319), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__3_ ( .D(
        mem_stage_inst_dmem_n1320), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__4_ ( .D(
        mem_stage_inst_dmem_n1321), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__5_ ( .D(
        mem_stage_inst_dmem_n1322), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__6_ ( .D(
        mem_stage_inst_dmem_n1323), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__7_ ( .D(
        mem_stage_inst_dmem_n1324), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__8_ ( .D(
        mem_stage_inst_dmem_n1325), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__9_ ( .D(
        mem_stage_inst_dmem_n1326), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__10_ ( .D(
        mem_stage_inst_dmem_n1327), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__11_ ( .D(
        mem_stage_inst_dmem_n1328), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__12_ ( .D(
        mem_stage_inst_dmem_n1329), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__13_ ( .D(
        mem_stage_inst_dmem_n1330), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__14_ ( .D(
        mem_stage_inst_dmem_n1331), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_47__15_ ( .D(
        mem_stage_inst_dmem_n1332), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_47__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__0_ ( .D(
        mem_stage_inst_dmem_n1381), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__1_ ( .D(
        mem_stage_inst_dmem_n1382), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__2_ ( .D(
        mem_stage_inst_dmem_n1383), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__3_ ( .D(
        mem_stage_inst_dmem_n1384), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__4_ ( .D(
        mem_stage_inst_dmem_n1385), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__5_ ( .D(
        mem_stage_inst_dmem_n1386), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__6_ ( .D(
        mem_stage_inst_dmem_n1387), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__7_ ( .D(
        mem_stage_inst_dmem_n1388), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__8_ ( .D(
        mem_stage_inst_dmem_n1389), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__9_ ( .D(
        mem_stage_inst_dmem_n1390), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__10_ ( .D(
        mem_stage_inst_dmem_n1391), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__11_ ( .D(
        mem_stage_inst_dmem_n1392), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__12_ ( .D(
        mem_stage_inst_dmem_n1393), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__13_ ( .D(
        mem_stage_inst_dmem_n1394), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__14_ ( .D(
        mem_stage_inst_dmem_n1395), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_51__15_ ( .D(
        mem_stage_inst_dmem_n1396), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_51__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__0_ ( .D(
        mem_stage_inst_dmem_n1445), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__1_ ( .D(
        mem_stage_inst_dmem_n1446), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__2_ ( .D(
        mem_stage_inst_dmem_n1447), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__3_ ( .D(
        mem_stage_inst_dmem_n1448), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__4_ ( .D(
        mem_stage_inst_dmem_n1449), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__5_ ( .D(
        mem_stage_inst_dmem_n1450), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__6_ ( .D(
        mem_stage_inst_dmem_n1451), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__7_ ( .D(
        mem_stage_inst_dmem_n1452), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__8_ ( .D(
        mem_stage_inst_dmem_n1453), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__9_ ( .D(
        mem_stage_inst_dmem_n1454), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__10_ ( .D(
        mem_stage_inst_dmem_n1455), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__11_ ( .D(
        mem_stage_inst_dmem_n1456), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__12_ ( .D(
        mem_stage_inst_dmem_n1457), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__13_ ( .D(
        mem_stage_inst_dmem_n1458), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__14_ ( .D(
        mem_stage_inst_dmem_n1459), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_55__15_ ( .D(
        mem_stage_inst_dmem_n1460), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_55__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__0_ ( .D(
        mem_stage_inst_dmem_n1509), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__1_ ( .D(
        mem_stage_inst_dmem_n1510), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__2_ ( .D(
        mem_stage_inst_dmem_n1511), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__3_ ( .D(
        mem_stage_inst_dmem_n1512), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__4_ ( .D(
        mem_stage_inst_dmem_n1513), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__5_ ( .D(
        mem_stage_inst_dmem_n1514), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__6_ ( .D(
        mem_stage_inst_dmem_n1515), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__7_ ( .D(
        mem_stage_inst_dmem_n1516), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__8_ ( .D(
        mem_stage_inst_dmem_n1517), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__9_ ( .D(
        mem_stage_inst_dmem_n1518), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__10_ ( .D(
        mem_stage_inst_dmem_n1519), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__11_ ( .D(
        mem_stage_inst_dmem_n1520), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__12_ ( .D(
        mem_stage_inst_dmem_n1521), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__13_ ( .D(
        mem_stage_inst_dmem_n1522), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__14_ ( .D(
        mem_stage_inst_dmem_n1523), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_59__15_ ( .D(
        mem_stage_inst_dmem_n1524), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_59__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__0_ ( .D(
        mem_stage_inst_dmem_n1573), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__1_ ( .D(
        mem_stage_inst_dmem_n1574), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__2_ ( .D(
        mem_stage_inst_dmem_n1575), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__3_ ( .D(
        mem_stage_inst_dmem_n1576), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__4_ ( .D(
        mem_stage_inst_dmem_n1577), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__5_ ( .D(
        mem_stage_inst_dmem_n1578), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__6_ ( .D(
        mem_stage_inst_dmem_n1579), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__7_ ( .D(
        mem_stage_inst_dmem_n1580), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__8_ ( .D(
        mem_stage_inst_dmem_n1581), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__9_ ( .D(
        mem_stage_inst_dmem_n1582), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__10_ ( .D(
        mem_stage_inst_dmem_n1583), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__11_ ( .D(
        mem_stage_inst_dmem_n1584), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__12_ ( .D(
        mem_stage_inst_dmem_n1585), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__13_ ( .D(
        mem_stage_inst_dmem_n1586), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__14_ ( .D(
        mem_stage_inst_dmem_n1587), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_63__15_ ( .D(
        mem_stage_inst_dmem_n1588), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_63__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__0_ ( .D(
        mem_stage_inst_dmem_n1637), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__1_ ( .D(
        mem_stage_inst_dmem_n1638), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__2_ ( .D(
        mem_stage_inst_dmem_n1639), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__3_ ( .D(
        mem_stage_inst_dmem_n1640), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__4_ ( .D(
        mem_stage_inst_dmem_n1641), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__5_ ( .D(
        mem_stage_inst_dmem_n1642), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__6_ ( .D(
        mem_stage_inst_dmem_n1643), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__7_ ( .D(
        mem_stage_inst_dmem_n1644), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__8_ ( .D(
        mem_stage_inst_dmem_n1645), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__9_ ( .D(
        mem_stage_inst_dmem_n1646), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__10_ ( .D(
        mem_stage_inst_dmem_n1647), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__11_ ( .D(
        mem_stage_inst_dmem_n1648), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__12_ ( .D(
        mem_stage_inst_dmem_n1649), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__13_ ( .D(
        mem_stage_inst_dmem_n1650), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__14_ ( .D(
        mem_stage_inst_dmem_n1651), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_67__15_ ( .D(
        mem_stage_inst_dmem_n1652), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_67__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__0_ ( .D(
        mem_stage_inst_dmem_n1701), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__1_ ( .D(
        mem_stage_inst_dmem_n1702), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__2_ ( .D(
        mem_stage_inst_dmem_n1703), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__3_ ( .D(
        mem_stage_inst_dmem_n1704), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__4_ ( .D(
        mem_stage_inst_dmem_n1705), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__5_ ( .D(
        mem_stage_inst_dmem_n1706), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__6_ ( .D(
        mem_stage_inst_dmem_n1707), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__7_ ( .D(
        mem_stage_inst_dmem_n1708), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__8_ ( .D(
        mem_stage_inst_dmem_n1709), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__9_ ( .D(
        mem_stage_inst_dmem_n1710), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__10_ ( .D(
        mem_stage_inst_dmem_n1711), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__11_ ( .D(
        mem_stage_inst_dmem_n1712), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__12_ ( .D(
        mem_stage_inst_dmem_n1713), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__13_ ( .D(
        mem_stage_inst_dmem_n1714), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__14_ ( .D(
        mem_stage_inst_dmem_n1715), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_71__15_ ( .D(
        mem_stage_inst_dmem_n1716), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_71__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__0_ ( .D(
        mem_stage_inst_dmem_n1765), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__1_ ( .D(
        mem_stage_inst_dmem_n1766), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__2_ ( .D(
        mem_stage_inst_dmem_n1767), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__3_ ( .D(
        mem_stage_inst_dmem_n1768), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__4_ ( .D(
        mem_stage_inst_dmem_n1769), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__5_ ( .D(
        mem_stage_inst_dmem_n1770), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__6_ ( .D(
        mem_stage_inst_dmem_n1771), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__7_ ( .D(
        mem_stage_inst_dmem_n1772), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__8_ ( .D(
        mem_stage_inst_dmem_n1773), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__9_ ( .D(
        mem_stage_inst_dmem_n1774), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__10_ ( .D(
        mem_stage_inst_dmem_n1775), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__11_ ( .D(
        mem_stage_inst_dmem_n1776), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__12_ ( .D(
        mem_stage_inst_dmem_n1777), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__13_ ( .D(
        mem_stage_inst_dmem_n1778), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__14_ ( .D(
        mem_stage_inst_dmem_n1779), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_75__15_ ( .D(
        mem_stage_inst_dmem_n1780), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_75__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__0_ ( .D(
        mem_stage_inst_dmem_n1829), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__1_ ( .D(
        mem_stage_inst_dmem_n1830), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__2_ ( .D(
        mem_stage_inst_dmem_n1831), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__3_ ( .D(
        mem_stage_inst_dmem_n1832), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__4_ ( .D(
        mem_stage_inst_dmem_n1833), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__5_ ( .D(
        mem_stage_inst_dmem_n1834), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__6_ ( .D(
        mem_stage_inst_dmem_n1835), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__7_ ( .D(
        mem_stage_inst_dmem_n1836), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__8_ ( .D(
        mem_stage_inst_dmem_n1837), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__9_ ( .D(
        mem_stage_inst_dmem_n1838), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__10_ ( .D(
        mem_stage_inst_dmem_n1839), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__11_ ( .D(
        mem_stage_inst_dmem_n1840), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__12_ ( .D(
        mem_stage_inst_dmem_n1841), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__13_ ( .D(
        mem_stage_inst_dmem_n1842), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__14_ ( .D(
        mem_stage_inst_dmem_n1843), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_79__15_ ( .D(
        mem_stage_inst_dmem_n1844), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_79__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__0_ ( .D(
        mem_stage_inst_dmem_n1893), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__1_ ( .D(
        mem_stage_inst_dmem_n1894), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__2_ ( .D(
        mem_stage_inst_dmem_n1895), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__3_ ( .D(
        mem_stage_inst_dmem_n1896), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__4_ ( .D(
        mem_stage_inst_dmem_n1897), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__5_ ( .D(
        mem_stage_inst_dmem_n1898), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__6_ ( .D(
        mem_stage_inst_dmem_n1899), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__7_ ( .D(
        mem_stage_inst_dmem_n1900), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__8_ ( .D(
        mem_stage_inst_dmem_n1901), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__9_ ( .D(
        mem_stage_inst_dmem_n1902), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__10_ ( .D(
        mem_stage_inst_dmem_n1903), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__11_ ( .D(
        mem_stage_inst_dmem_n1904), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__12_ ( .D(
        mem_stage_inst_dmem_n1905), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__13_ ( .D(
        mem_stage_inst_dmem_n1906), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__14_ ( .D(
        mem_stage_inst_dmem_n1907), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_83__15_ ( .D(
        mem_stage_inst_dmem_n1908), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_83__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__0_ ( .D(
        mem_stage_inst_dmem_n1957), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__1_ ( .D(
        mem_stage_inst_dmem_n1958), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__2_ ( .D(
        mem_stage_inst_dmem_n1959), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__3_ ( .D(
        mem_stage_inst_dmem_n1960), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__4_ ( .D(
        mem_stage_inst_dmem_n1961), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__5_ ( .D(
        mem_stage_inst_dmem_n1962), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__6_ ( .D(
        mem_stage_inst_dmem_n1963), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__7_ ( .D(
        mem_stage_inst_dmem_n1964), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__8_ ( .D(
        mem_stage_inst_dmem_n1965), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__9_ ( .D(
        mem_stage_inst_dmem_n1966), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__10_ ( .D(
        mem_stage_inst_dmem_n1967), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__11_ ( .D(
        mem_stage_inst_dmem_n1968), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__12_ ( .D(
        mem_stage_inst_dmem_n1969), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__13_ ( .D(
        mem_stage_inst_dmem_n1970), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__14_ ( .D(
        mem_stage_inst_dmem_n1971), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_87__15_ ( .D(
        mem_stage_inst_dmem_n1972), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_87__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__0_ ( .D(
        mem_stage_inst_dmem_n2021), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__1_ ( .D(
        mem_stage_inst_dmem_n2022), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__2_ ( .D(
        mem_stage_inst_dmem_n2023), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__3_ ( .D(
        mem_stage_inst_dmem_n2024), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__4_ ( .D(
        mem_stage_inst_dmem_n2025), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__5_ ( .D(
        mem_stage_inst_dmem_n2026), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__6_ ( .D(
        mem_stage_inst_dmem_n2027), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__7_ ( .D(
        mem_stage_inst_dmem_n2028), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__8_ ( .D(
        mem_stage_inst_dmem_n2029), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__9_ ( .D(
        mem_stage_inst_dmem_n2030), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__10_ ( .D(
        mem_stage_inst_dmem_n2031), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__11_ ( .D(
        mem_stage_inst_dmem_n2032), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__12_ ( .D(
        mem_stage_inst_dmem_n2033), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__13_ ( .D(
        mem_stage_inst_dmem_n2034), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__14_ ( .D(
        mem_stage_inst_dmem_n2035), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_91__15_ ( .D(
        mem_stage_inst_dmem_n2036), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_91__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__0_ ( .D(
        mem_stage_inst_dmem_n2085), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__1_ ( .D(
        mem_stage_inst_dmem_n2086), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__2_ ( .D(
        mem_stage_inst_dmem_n2087), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__3_ ( .D(
        mem_stage_inst_dmem_n2088), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__4_ ( .D(
        mem_stage_inst_dmem_n2089), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__5_ ( .D(
        mem_stage_inst_dmem_n2090), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__6_ ( .D(
        mem_stage_inst_dmem_n2091), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__7_ ( .D(
        mem_stage_inst_dmem_n2092), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__8_ ( .D(
        mem_stage_inst_dmem_n2093), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__9_ ( .D(
        mem_stage_inst_dmem_n2094), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__10_ ( .D(
        mem_stage_inst_dmem_n2095), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__11_ ( .D(
        mem_stage_inst_dmem_n2096), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__12_ ( .D(
        mem_stage_inst_dmem_n2097), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__13_ ( .D(
        mem_stage_inst_dmem_n2098), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__14_ ( .D(
        mem_stage_inst_dmem_n2099), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_95__15_ ( .D(
        mem_stage_inst_dmem_n2100), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_95__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__0_ ( .D(
        mem_stage_inst_dmem_n2149), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__1_ ( .D(
        mem_stage_inst_dmem_n2150), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__2_ ( .D(
        mem_stage_inst_dmem_n2151), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__3_ ( .D(
        mem_stage_inst_dmem_n2152), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__4_ ( .D(
        mem_stage_inst_dmem_n2153), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__5_ ( .D(
        mem_stage_inst_dmem_n2154), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__6_ ( .D(
        mem_stage_inst_dmem_n2155), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__7_ ( .D(
        mem_stage_inst_dmem_n2156), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__8_ ( .D(
        mem_stage_inst_dmem_n2157), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__9_ ( .D(
        mem_stage_inst_dmem_n2158), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__10_ ( .D(
        mem_stage_inst_dmem_n2159), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__11_ ( .D(
        mem_stage_inst_dmem_n2160), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__12_ ( .D(
        mem_stage_inst_dmem_n2161), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__13_ ( .D(
        mem_stage_inst_dmem_n2162), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__14_ ( .D(
        mem_stage_inst_dmem_n2163), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_99__15_ ( .D(
        mem_stage_inst_dmem_n2164), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_99__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__0_ ( .D(
        mem_stage_inst_dmem_n2213), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__1_ ( .D(
        mem_stage_inst_dmem_n2214), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__2_ ( .D(
        mem_stage_inst_dmem_n2215), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__3_ ( .D(
        mem_stage_inst_dmem_n2216), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__4_ ( .D(
        mem_stage_inst_dmem_n2217), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__5_ ( .D(
        mem_stage_inst_dmem_n2218), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__6_ ( .D(
        mem_stage_inst_dmem_n2219), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__7_ ( .D(
        mem_stage_inst_dmem_n2220), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__8_ ( .D(
        mem_stage_inst_dmem_n2221), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__9_ ( .D(
        mem_stage_inst_dmem_n2222), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__10_ ( .D(
        mem_stage_inst_dmem_n2223), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__11_ ( .D(
        mem_stage_inst_dmem_n2224), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__12_ ( .D(
        mem_stage_inst_dmem_n2225), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__13_ ( .D(
        mem_stage_inst_dmem_n2226), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__14_ ( .D(
        mem_stage_inst_dmem_n2227), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_103__15_ ( .D(
        mem_stage_inst_dmem_n2228), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_103__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__0_ ( .D(
        mem_stage_inst_dmem_n2277), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__1_ ( .D(
        mem_stage_inst_dmem_n2278), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__2_ ( .D(
        mem_stage_inst_dmem_n2279), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__3_ ( .D(
        mem_stage_inst_dmem_n2280), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__4_ ( .D(
        mem_stage_inst_dmem_n2281), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__5_ ( .D(
        mem_stage_inst_dmem_n2282), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__6_ ( .D(
        mem_stage_inst_dmem_n2283), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__7_ ( .D(
        mem_stage_inst_dmem_n2284), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__8_ ( .D(
        mem_stage_inst_dmem_n2285), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__9_ ( .D(
        mem_stage_inst_dmem_n2286), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__10_ ( .D(
        mem_stage_inst_dmem_n2287), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__11_ ( .D(
        mem_stage_inst_dmem_n2288), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__12_ ( .D(
        mem_stage_inst_dmem_n2289), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__13_ ( .D(
        mem_stage_inst_dmem_n2290), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__14_ ( .D(
        mem_stage_inst_dmem_n2291), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_107__15_ ( .D(
        mem_stage_inst_dmem_n2292), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_107__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__0_ ( .D(
        mem_stage_inst_dmem_n2341), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__1_ ( .D(
        mem_stage_inst_dmem_n2342), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__2_ ( .D(
        mem_stage_inst_dmem_n2343), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__3_ ( .D(
        mem_stage_inst_dmem_n2344), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__4_ ( .D(
        mem_stage_inst_dmem_n2345), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__5_ ( .D(
        mem_stage_inst_dmem_n2346), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__6_ ( .D(
        mem_stage_inst_dmem_n2347), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__7_ ( .D(
        mem_stage_inst_dmem_n2348), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__8_ ( .D(
        mem_stage_inst_dmem_n2349), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__9_ ( .D(
        mem_stage_inst_dmem_n2350), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__10_ ( .D(
        mem_stage_inst_dmem_n2351), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__11_ ( .D(
        mem_stage_inst_dmem_n2352), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__12_ ( .D(
        mem_stage_inst_dmem_n2353), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__13_ ( .D(
        mem_stage_inst_dmem_n2354), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__14_ ( .D(
        mem_stage_inst_dmem_n2355), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_111__15_ ( .D(
        mem_stage_inst_dmem_n2356), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_111__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__0_ ( .D(
        mem_stage_inst_dmem_n2405), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__1_ ( .D(
        mem_stage_inst_dmem_n2406), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__2_ ( .D(
        mem_stage_inst_dmem_n2407), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__3_ ( .D(
        mem_stage_inst_dmem_n2408), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__4_ ( .D(
        mem_stage_inst_dmem_n2409), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__5_ ( .D(
        mem_stage_inst_dmem_n2410), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__6_ ( .D(
        mem_stage_inst_dmem_n2411), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__7_ ( .D(
        mem_stage_inst_dmem_n2412), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__8_ ( .D(
        mem_stage_inst_dmem_n2413), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__9_ ( .D(
        mem_stage_inst_dmem_n2414), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__10_ ( .D(
        mem_stage_inst_dmem_n2415), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__11_ ( .D(
        mem_stage_inst_dmem_n2416), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__12_ ( .D(
        mem_stage_inst_dmem_n2417), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__13_ ( .D(
        mem_stage_inst_dmem_n2418), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__14_ ( .D(
        mem_stage_inst_dmem_n2419), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_115__15_ ( .D(
        mem_stage_inst_dmem_n2420), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_115__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__0_ ( .D(
        mem_stage_inst_dmem_n2469), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__1_ ( .D(
        mem_stage_inst_dmem_n2470), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__2_ ( .D(
        mem_stage_inst_dmem_n2471), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__3_ ( .D(
        mem_stage_inst_dmem_n2472), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__4_ ( .D(
        mem_stage_inst_dmem_n2473), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__5_ ( .D(
        mem_stage_inst_dmem_n2474), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__6_ ( .D(
        mem_stage_inst_dmem_n2475), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__7_ ( .D(
        mem_stage_inst_dmem_n2476), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__8_ ( .D(
        mem_stage_inst_dmem_n2477), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__9_ ( .D(
        mem_stage_inst_dmem_n2478), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__10_ ( .D(
        mem_stage_inst_dmem_n2479), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__11_ ( .D(
        mem_stage_inst_dmem_n2480), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__12_ ( .D(
        mem_stage_inst_dmem_n2481), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__13_ ( .D(
        mem_stage_inst_dmem_n2482), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__14_ ( .D(
        mem_stage_inst_dmem_n2483), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_119__15_ ( .D(
        mem_stage_inst_dmem_n2484), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_119__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__0_ ( .D(
        mem_stage_inst_dmem_n2533), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__1_ ( .D(
        mem_stage_inst_dmem_n2534), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__2_ ( .D(
        mem_stage_inst_dmem_n2535), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__3_ ( .D(
        mem_stage_inst_dmem_n2536), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__4_ ( .D(
        mem_stage_inst_dmem_n2537), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__5_ ( .D(
        mem_stage_inst_dmem_n2538), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__6_ ( .D(
        mem_stage_inst_dmem_n2539), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__7_ ( .D(
        mem_stage_inst_dmem_n2540), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__8_ ( .D(
        mem_stage_inst_dmem_n2541), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__9_ ( .D(
        mem_stage_inst_dmem_n2542), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__10_ ( .D(
        mem_stage_inst_dmem_n2543), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__11_ ( .D(
        mem_stage_inst_dmem_n2544), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__12_ ( .D(
        mem_stage_inst_dmem_n2545), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__13_ ( .D(
        mem_stage_inst_dmem_n2546), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__14_ ( .D(
        mem_stage_inst_dmem_n2547), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_123__15_ ( .D(
        mem_stage_inst_dmem_n2548), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_123__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__0_ ( .D(
        mem_stage_inst_dmem_n2597), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__1_ ( .D(
        mem_stage_inst_dmem_n2598), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__2_ ( .D(
        mem_stage_inst_dmem_n2599), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__3_ ( .D(
        mem_stage_inst_dmem_n2600), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__4_ ( .D(
        mem_stage_inst_dmem_n2601), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__5_ ( .D(
        mem_stage_inst_dmem_n2602), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__6_ ( .D(
        mem_stage_inst_dmem_n2603), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__7_ ( .D(
        mem_stage_inst_dmem_n2604), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__8_ ( .D(
        mem_stage_inst_dmem_n2605), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__9_ ( .D(
        mem_stage_inst_dmem_n2606), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__10_ ( .D(
        mem_stage_inst_dmem_n2607), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__11_ ( .D(
        mem_stage_inst_dmem_n2608), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__12_ ( .D(
        mem_stage_inst_dmem_n2609), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__13_ ( .D(
        mem_stage_inst_dmem_n2610), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__14_ ( .D(
        mem_stage_inst_dmem_n2611), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_127__15_ ( .D(
        mem_stage_inst_dmem_n2612), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_127__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__0_ ( .D(
        mem_stage_inst_dmem_n2661), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__1_ ( .D(
        mem_stage_inst_dmem_n2662), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__2_ ( .D(
        mem_stage_inst_dmem_n2663), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__3_ ( .D(
        mem_stage_inst_dmem_n2664), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__4_ ( .D(
        mem_stage_inst_dmem_n2665), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__5_ ( .D(
        mem_stage_inst_dmem_n2666), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__6_ ( .D(
        mem_stage_inst_dmem_n2667), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__7_ ( .D(
        mem_stage_inst_dmem_n2668), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__8_ ( .D(
        mem_stage_inst_dmem_n2669), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__9_ ( .D(
        mem_stage_inst_dmem_n2670), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__10_ ( .D(
        mem_stage_inst_dmem_n2671), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__11_ ( .D(
        mem_stage_inst_dmem_n2672), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__12_ ( .D(
        mem_stage_inst_dmem_n2673), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__13_ ( .D(
        mem_stage_inst_dmem_n2674), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__14_ ( .D(
        mem_stage_inst_dmem_n2675), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_131__15_ ( .D(
        mem_stage_inst_dmem_n2676), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_131__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__0_ ( .D(
        mem_stage_inst_dmem_n2725), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__1_ ( .D(
        mem_stage_inst_dmem_n2726), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__2_ ( .D(
        mem_stage_inst_dmem_n2727), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__3_ ( .D(
        mem_stage_inst_dmem_n2728), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__4_ ( .D(
        mem_stage_inst_dmem_n2729), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__5_ ( .D(
        mem_stage_inst_dmem_n2730), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__6_ ( .D(
        mem_stage_inst_dmem_n2731), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__7_ ( .D(
        mem_stage_inst_dmem_n2732), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__8_ ( .D(
        mem_stage_inst_dmem_n2733), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__9_ ( .D(
        mem_stage_inst_dmem_n2734), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__10_ ( .D(
        mem_stage_inst_dmem_n2735), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__11_ ( .D(
        mem_stage_inst_dmem_n2736), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__12_ ( .D(
        mem_stage_inst_dmem_n2737), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__13_ ( .D(
        mem_stage_inst_dmem_n2738), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__14_ ( .D(
        mem_stage_inst_dmem_n2739), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_135__15_ ( .D(
        mem_stage_inst_dmem_n2740), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_135__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__0_ ( .D(
        mem_stage_inst_dmem_n2789), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__1_ ( .D(
        mem_stage_inst_dmem_n2790), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__2_ ( .D(
        mem_stage_inst_dmem_n2791), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__3_ ( .D(
        mem_stage_inst_dmem_n2792), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__4_ ( .D(
        mem_stage_inst_dmem_n2793), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__5_ ( .D(
        mem_stage_inst_dmem_n2794), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__6_ ( .D(
        mem_stage_inst_dmem_n2795), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__7_ ( .D(
        mem_stage_inst_dmem_n2796), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__8_ ( .D(
        mem_stage_inst_dmem_n2797), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__9_ ( .D(
        mem_stage_inst_dmem_n2798), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__10_ ( .D(
        mem_stage_inst_dmem_n2799), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__11_ ( .D(
        mem_stage_inst_dmem_n2800), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__12_ ( .D(
        mem_stage_inst_dmem_n2801), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__13_ ( .D(
        mem_stage_inst_dmem_n2802), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__14_ ( .D(
        mem_stage_inst_dmem_n2803), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_139__15_ ( .D(
        mem_stage_inst_dmem_n2804), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_139__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__0_ ( .D(
        mem_stage_inst_dmem_n2853), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__1_ ( .D(
        mem_stage_inst_dmem_n2854), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__2_ ( .D(
        mem_stage_inst_dmem_n2855), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__3_ ( .D(
        mem_stage_inst_dmem_n2856), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__4_ ( .D(
        mem_stage_inst_dmem_n2857), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__5_ ( .D(
        mem_stage_inst_dmem_n2858), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__6_ ( .D(
        mem_stage_inst_dmem_n2859), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__7_ ( .D(
        mem_stage_inst_dmem_n2860), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__8_ ( .D(
        mem_stage_inst_dmem_n2861), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__9_ ( .D(
        mem_stage_inst_dmem_n2862), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__10_ ( .D(
        mem_stage_inst_dmem_n2863), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__11_ ( .D(
        mem_stage_inst_dmem_n2864), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__12_ ( .D(
        mem_stage_inst_dmem_n2865), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__13_ ( .D(
        mem_stage_inst_dmem_n2866), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__14_ ( .D(
        mem_stage_inst_dmem_n2867), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_143__15_ ( .D(
        mem_stage_inst_dmem_n2868), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_143__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__0_ ( .D(
        mem_stage_inst_dmem_n2917), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__1_ ( .D(
        mem_stage_inst_dmem_n2918), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__2_ ( .D(
        mem_stage_inst_dmem_n2919), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__3_ ( .D(
        mem_stage_inst_dmem_n2920), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__4_ ( .D(
        mem_stage_inst_dmem_n2921), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__5_ ( .D(
        mem_stage_inst_dmem_n2922), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__6_ ( .D(
        mem_stage_inst_dmem_n2923), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__7_ ( .D(
        mem_stage_inst_dmem_n2924), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__8_ ( .D(
        mem_stage_inst_dmem_n2925), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__9_ ( .D(
        mem_stage_inst_dmem_n2926), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__10_ ( .D(
        mem_stage_inst_dmem_n2927), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__11_ ( .D(
        mem_stage_inst_dmem_n2928), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__12_ ( .D(
        mem_stage_inst_dmem_n2929), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__13_ ( .D(
        mem_stage_inst_dmem_n2930), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__14_ ( .D(
        mem_stage_inst_dmem_n2931), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_147__15_ ( .D(
        mem_stage_inst_dmem_n2932), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_147__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__0_ ( .D(
        mem_stage_inst_dmem_n2981), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__1_ ( .D(
        mem_stage_inst_dmem_n2982), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__2_ ( .D(
        mem_stage_inst_dmem_n2983), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__3_ ( .D(
        mem_stage_inst_dmem_n2984), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__4_ ( .D(
        mem_stage_inst_dmem_n2985), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__5_ ( .D(
        mem_stage_inst_dmem_n2986), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__6_ ( .D(
        mem_stage_inst_dmem_n2987), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__7_ ( .D(
        mem_stage_inst_dmem_n2988), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__8_ ( .D(
        mem_stage_inst_dmem_n2989), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__9_ ( .D(
        mem_stage_inst_dmem_n2990), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__10_ ( .D(
        mem_stage_inst_dmem_n2991), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__11_ ( .D(
        mem_stage_inst_dmem_n2992), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__12_ ( .D(
        mem_stage_inst_dmem_n2993), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__13_ ( .D(
        mem_stage_inst_dmem_n2994), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__14_ ( .D(
        mem_stage_inst_dmem_n2995), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_151__15_ ( .D(
        mem_stage_inst_dmem_n2996), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_151__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__0_ ( .D(
        mem_stage_inst_dmem_n3045), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__1_ ( .D(
        mem_stage_inst_dmem_n3046), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__2_ ( .D(
        mem_stage_inst_dmem_n3047), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__3_ ( .D(
        mem_stage_inst_dmem_n3048), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__4_ ( .D(
        mem_stage_inst_dmem_n3049), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__5_ ( .D(
        mem_stage_inst_dmem_n3050), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__6_ ( .D(
        mem_stage_inst_dmem_n3051), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__7_ ( .D(
        mem_stage_inst_dmem_n3052), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__8_ ( .D(
        mem_stage_inst_dmem_n3053), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__9_ ( .D(
        mem_stage_inst_dmem_n3054), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__10_ ( .D(
        mem_stage_inst_dmem_n3055), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__11_ ( .D(
        mem_stage_inst_dmem_n3056), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__12_ ( .D(
        mem_stage_inst_dmem_n3057), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__13_ ( .D(
        mem_stage_inst_dmem_n3058), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__14_ ( .D(
        mem_stage_inst_dmem_n3059), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_155__15_ ( .D(
        mem_stage_inst_dmem_n3060), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_155__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__0_ ( .D(
        mem_stage_inst_dmem_n3109), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__1_ ( .D(
        mem_stage_inst_dmem_n3110), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__2_ ( .D(
        mem_stage_inst_dmem_n3111), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__3_ ( .D(
        mem_stage_inst_dmem_n3112), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__4_ ( .D(
        mem_stage_inst_dmem_n3113), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__5_ ( .D(
        mem_stage_inst_dmem_n3114), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__6_ ( .D(
        mem_stage_inst_dmem_n3115), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__7_ ( .D(
        mem_stage_inst_dmem_n3116), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__8_ ( .D(
        mem_stage_inst_dmem_n3117), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__9_ ( .D(
        mem_stage_inst_dmem_n3118), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__10_ ( .D(
        mem_stage_inst_dmem_n3119), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__11_ ( .D(
        mem_stage_inst_dmem_n3120), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__12_ ( .D(
        mem_stage_inst_dmem_n3121), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__13_ ( .D(
        mem_stage_inst_dmem_n3122), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__14_ ( .D(
        mem_stage_inst_dmem_n3123), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_159__15_ ( .D(
        mem_stage_inst_dmem_n3124), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_159__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__0_ ( .D(
        mem_stage_inst_dmem_n3173), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__1_ ( .D(
        mem_stage_inst_dmem_n3174), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__2_ ( .D(
        mem_stage_inst_dmem_n3175), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__3_ ( .D(
        mem_stage_inst_dmem_n3176), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__4_ ( .D(
        mem_stage_inst_dmem_n3177), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__5_ ( .D(
        mem_stage_inst_dmem_n3178), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__6_ ( .D(
        mem_stage_inst_dmem_n3179), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__7_ ( .D(
        mem_stage_inst_dmem_n3180), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__8_ ( .D(
        mem_stage_inst_dmem_n3181), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__9_ ( .D(
        mem_stage_inst_dmem_n3182), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__10_ ( .D(
        mem_stage_inst_dmem_n3183), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__11_ ( .D(
        mem_stage_inst_dmem_n3184), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__12_ ( .D(
        mem_stage_inst_dmem_n3185), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__13_ ( .D(
        mem_stage_inst_dmem_n3186), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__14_ ( .D(
        mem_stage_inst_dmem_n3187), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_163__15_ ( .D(
        mem_stage_inst_dmem_n3188), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_163__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__0_ ( .D(
        mem_stage_inst_dmem_n3237), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__1_ ( .D(
        mem_stage_inst_dmem_n3238), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__2_ ( .D(
        mem_stage_inst_dmem_n3239), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__3_ ( .D(
        mem_stage_inst_dmem_n3240), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__4_ ( .D(
        mem_stage_inst_dmem_n3241), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__5_ ( .D(
        mem_stage_inst_dmem_n3242), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__6_ ( .D(
        mem_stage_inst_dmem_n3243), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__7_ ( .D(
        mem_stage_inst_dmem_n3244), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__8_ ( .D(
        mem_stage_inst_dmem_n3245), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__9_ ( .D(
        mem_stage_inst_dmem_n3246), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__10_ ( .D(
        mem_stage_inst_dmem_n3247), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__11_ ( .D(
        mem_stage_inst_dmem_n3248), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__12_ ( .D(
        mem_stage_inst_dmem_n3249), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__13_ ( .D(
        mem_stage_inst_dmem_n3250), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__14_ ( .D(
        mem_stage_inst_dmem_n3251), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_167__15_ ( .D(
        mem_stage_inst_dmem_n3252), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_167__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__0_ ( .D(
        mem_stage_inst_dmem_n3301), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__1_ ( .D(
        mem_stage_inst_dmem_n3302), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__2_ ( .D(
        mem_stage_inst_dmem_n3303), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__3_ ( .D(
        mem_stage_inst_dmem_n3304), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__4_ ( .D(
        mem_stage_inst_dmem_n3305), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__5_ ( .D(
        mem_stage_inst_dmem_n3306), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__6_ ( .D(
        mem_stage_inst_dmem_n3307), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__7_ ( .D(
        mem_stage_inst_dmem_n3308), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__8_ ( .D(
        mem_stage_inst_dmem_n3309), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__9_ ( .D(
        mem_stage_inst_dmem_n3310), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__10_ ( .D(
        mem_stage_inst_dmem_n3311), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__11_ ( .D(
        mem_stage_inst_dmem_n3312), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__12_ ( .D(
        mem_stage_inst_dmem_n3313), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__13_ ( .D(
        mem_stage_inst_dmem_n3314), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__14_ ( .D(
        mem_stage_inst_dmem_n3315), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_171__15_ ( .D(
        mem_stage_inst_dmem_n3316), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_171__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__0_ ( .D(
        mem_stage_inst_dmem_n3365), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__1_ ( .D(
        mem_stage_inst_dmem_n3366), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__2_ ( .D(
        mem_stage_inst_dmem_n3367), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__3_ ( .D(
        mem_stage_inst_dmem_n3368), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__4_ ( .D(
        mem_stage_inst_dmem_n3369), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__5_ ( .D(
        mem_stage_inst_dmem_n3370), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__6_ ( .D(
        mem_stage_inst_dmem_n3371), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__7_ ( .D(
        mem_stage_inst_dmem_n3372), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__8_ ( .D(
        mem_stage_inst_dmem_n3373), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__9_ ( .D(
        mem_stage_inst_dmem_n3374), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__10_ ( .D(
        mem_stage_inst_dmem_n3375), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__11_ ( .D(
        mem_stage_inst_dmem_n3376), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__12_ ( .D(
        mem_stage_inst_dmem_n3377), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__13_ ( .D(
        mem_stage_inst_dmem_n3378), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__14_ ( .D(
        mem_stage_inst_dmem_n3379), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_175__15_ ( .D(
        mem_stage_inst_dmem_n3380), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_175__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__0_ ( .D(
        mem_stage_inst_dmem_n3429), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__1_ ( .D(
        mem_stage_inst_dmem_n3430), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__2_ ( .D(
        mem_stage_inst_dmem_n3431), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__3_ ( .D(
        mem_stage_inst_dmem_n3432), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__4_ ( .D(
        mem_stage_inst_dmem_n3433), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__5_ ( .D(
        mem_stage_inst_dmem_n3434), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__6_ ( .D(
        mem_stage_inst_dmem_n3435), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__7_ ( .D(
        mem_stage_inst_dmem_n3436), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__8_ ( .D(
        mem_stage_inst_dmem_n3437), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__9_ ( .D(
        mem_stage_inst_dmem_n3438), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__10_ ( .D(
        mem_stage_inst_dmem_n3439), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__11_ ( .D(
        mem_stage_inst_dmem_n3440), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__12_ ( .D(
        mem_stage_inst_dmem_n3441), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__13_ ( .D(
        mem_stage_inst_dmem_n3442), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__14_ ( .D(
        mem_stage_inst_dmem_n3443), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_179__15_ ( .D(
        mem_stage_inst_dmem_n3444), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_179__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__0_ ( .D(
        mem_stage_inst_dmem_n3493), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__1_ ( .D(
        mem_stage_inst_dmem_n3494), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__2_ ( .D(
        mem_stage_inst_dmem_n3495), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__3_ ( .D(
        mem_stage_inst_dmem_n3496), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__4_ ( .D(
        mem_stage_inst_dmem_n3497), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__5_ ( .D(
        mem_stage_inst_dmem_n3498), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__6_ ( .D(
        mem_stage_inst_dmem_n3499), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__7_ ( .D(
        mem_stage_inst_dmem_n3500), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__8_ ( .D(
        mem_stage_inst_dmem_n3501), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__9_ ( .D(
        mem_stage_inst_dmem_n3502), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__10_ ( .D(
        mem_stage_inst_dmem_n3503), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__11_ ( .D(
        mem_stage_inst_dmem_n3504), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__12_ ( .D(
        mem_stage_inst_dmem_n3505), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__13_ ( .D(
        mem_stage_inst_dmem_n3506), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__14_ ( .D(
        mem_stage_inst_dmem_n3507), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_183__15_ ( .D(
        mem_stage_inst_dmem_n3508), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_183__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__0_ ( .D(
        mem_stage_inst_dmem_n3557), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__1_ ( .D(
        mem_stage_inst_dmem_n3558), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__2_ ( .D(
        mem_stage_inst_dmem_n3559), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__3_ ( .D(
        mem_stage_inst_dmem_n3560), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__4_ ( .D(
        mem_stage_inst_dmem_n3561), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__5_ ( .D(
        mem_stage_inst_dmem_n3562), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__6_ ( .D(
        mem_stage_inst_dmem_n3563), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__7_ ( .D(
        mem_stage_inst_dmem_n3564), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__8_ ( .D(
        mem_stage_inst_dmem_n3565), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__9_ ( .D(
        mem_stage_inst_dmem_n3566), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__10_ ( .D(
        mem_stage_inst_dmem_n3567), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__11_ ( .D(
        mem_stage_inst_dmem_n3568), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__12_ ( .D(
        mem_stage_inst_dmem_n3569), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__13_ ( .D(
        mem_stage_inst_dmem_n3570), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__14_ ( .D(
        mem_stage_inst_dmem_n3571), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_187__15_ ( .D(
        mem_stage_inst_dmem_n3572), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_187__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__0_ ( .D(
        mem_stage_inst_dmem_n3621), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__1_ ( .D(
        mem_stage_inst_dmem_n3622), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__2_ ( .D(
        mem_stage_inst_dmem_n3623), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__3_ ( .D(
        mem_stage_inst_dmem_n3624), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__4_ ( .D(
        mem_stage_inst_dmem_n3625), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__5_ ( .D(
        mem_stage_inst_dmem_n3626), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__6_ ( .D(
        mem_stage_inst_dmem_n3627), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__7_ ( .D(
        mem_stage_inst_dmem_n3628), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__8_ ( .D(
        mem_stage_inst_dmem_n3629), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__9_ ( .D(
        mem_stage_inst_dmem_n3630), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__10_ ( .D(
        mem_stage_inst_dmem_n3631), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__11_ ( .D(
        mem_stage_inst_dmem_n3632), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__12_ ( .D(
        mem_stage_inst_dmem_n3633), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__13_ ( .D(
        mem_stage_inst_dmem_n3634), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__14_ ( .D(
        mem_stage_inst_dmem_n3635), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_191__15_ ( .D(
        mem_stage_inst_dmem_n3636), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_191__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__0_ ( .D(
        mem_stage_inst_dmem_n3685), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__1_ ( .D(
        mem_stage_inst_dmem_n3686), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__2_ ( .D(
        mem_stage_inst_dmem_n3687), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__3_ ( .D(
        mem_stage_inst_dmem_n3688), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__4_ ( .D(
        mem_stage_inst_dmem_n3689), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__5_ ( .D(
        mem_stage_inst_dmem_n3690), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__6_ ( .D(
        mem_stage_inst_dmem_n3691), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__7_ ( .D(
        mem_stage_inst_dmem_n3692), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__8_ ( .D(
        mem_stage_inst_dmem_n3693), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__9_ ( .D(
        mem_stage_inst_dmem_n3694), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__10_ ( .D(
        mem_stage_inst_dmem_n3695), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__11_ ( .D(
        mem_stage_inst_dmem_n3696), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__12_ ( .D(
        mem_stage_inst_dmem_n3697), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__13_ ( .D(
        mem_stage_inst_dmem_n3698), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__14_ ( .D(
        mem_stage_inst_dmem_n3699), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_195__15_ ( .D(
        mem_stage_inst_dmem_n3700), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_195__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__0_ ( .D(
        mem_stage_inst_dmem_n3749), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__1_ ( .D(
        mem_stage_inst_dmem_n3750), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__2_ ( .D(
        mem_stage_inst_dmem_n3751), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__3_ ( .D(
        mem_stage_inst_dmem_n3752), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__4_ ( .D(
        mem_stage_inst_dmem_n3753), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__5_ ( .D(
        mem_stage_inst_dmem_n3754), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__6_ ( .D(
        mem_stage_inst_dmem_n3755), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__7_ ( .D(
        mem_stage_inst_dmem_n3756), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__8_ ( .D(
        mem_stage_inst_dmem_n3757), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__9_ ( .D(
        mem_stage_inst_dmem_n3758), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__10_ ( .D(
        mem_stage_inst_dmem_n3759), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__11_ ( .D(
        mem_stage_inst_dmem_n3760), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__12_ ( .D(
        mem_stage_inst_dmem_n3761), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__13_ ( .D(
        mem_stage_inst_dmem_n3762), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__14_ ( .D(
        mem_stage_inst_dmem_n3763), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_199__15_ ( .D(
        mem_stage_inst_dmem_n3764), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_199__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__0_ ( .D(
        mem_stage_inst_dmem_n3813), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__1_ ( .D(
        mem_stage_inst_dmem_n3814), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__2_ ( .D(
        mem_stage_inst_dmem_n3815), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__3_ ( .D(
        mem_stage_inst_dmem_n3816), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__4_ ( .D(
        mem_stage_inst_dmem_n3817), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__5_ ( .D(
        mem_stage_inst_dmem_n3818), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__6_ ( .D(
        mem_stage_inst_dmem_n3819), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__7_ ( .D(
        mem_stage_inst_dmem_n3820), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__8_ ( .D(
        mem_stage_inst_dmem_n3821), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__9_ ( .D(
        mem_stage_inst_dmem_n3822), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__10_ ( .D(
        mem_stage_inst_dmem_n3823), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__11_ ( .D(
        mem_stage_inst_dmem_n3824), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__12_ ( .D(
        mem_stage_inst_dmem_n3825), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__13_ ( .D(
        mem_stage_inst_dmem_n3826), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__14_ ( .D(
        mem_stage_inst_dmem_n3827), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_203__15_ ( .D(
        mem_stage_inst_dmem_n3828), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_203__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__0_ ( .D(
        mem_stage_inst_dmem_n3877), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__1_ ( .D(
        mem_stage_inst_dmem_n3878), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__2_ ( .D(
        mem_stage_inst_dmem_n3879), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__3_ ( .D(
        mem_stage_inst_dmem_n3880), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__4_ ( .D(
        mem_stage_inst_dmem_n3881), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__5_ ( .D(
        mem_stage_inst_dmem_n3882), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__6_ ( .D(
        mem_stage_inst_dmem_n3883), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__7_ ( .D(
        mem_stage_inst_dmem_n3884), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__8_ ( .D(
        mem_stage_inst_dmem_n3885), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__9_ ( .D(
        mem_stage_inst_dmem_n3886), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__10_ ( .D(
        mem_stage_inst_dmem_n3887), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__11_ ( .D(
        mem_stage_inst_dmem_n3888), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__12_ ( .D(
        mem_stage_inst_dmem_n3889), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__13_ ( .D(
        mem_stage_inst_dmem_n3890), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__14_ ( .D(
        mem_stage_inst_dmem_n3891), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_207__15_ ( .D(
        mem_stage_inst_dmem_n3892), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_207__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__0_ ( .D(
        mem_stage_inst_dmem_n3941), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__1_ ( .D(
        mem_stage_inst_dmem_n3942), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__2_ ( .D(
        mem_stage_inst_dmem_n3943), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__3_ ( .D(
        mem_stage_inst_dmem_n3944), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__4_ ( .D(
        mem_stage_inst_dmem_n3945), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__5_ ( .D(
        mem_stage_inst_dmem_n3946), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__6_ ( .D(
        mem_stage_inst_dmem_n3947), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__7_ ( .D(
        mem_stage_inst_dmem_n3948), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__8_ ( .D(
        mem_stage_inst_dmem_n3949), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__9_ ( .D(
        mem_stage_inst_dmem_n3950), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__10_ ( .D(
        mem_stage_inst_dmem_n3951), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__11_ ( .D(
        mem_stage_inst_dmem_n3952), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__12_ ( .D(
        mem_stage_inst_dmem_n3953), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__13_ ( .D(
        mem_stage_inst_dmem_n3954), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__14_ ( .D(
        mem_stage_inst_dmem_n3955), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_211__15_ ( .D(
        mem_stage_inst_dmem_n3956), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_211__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__0_ ( .D(
        mem_stage_inst_dmem_n4005), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__1_ ( .D(
        mem_stage_inst_dmem_n4006), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__2_ ( .D(
        mem_stage_inst_dmem_n4007), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__3_ ( .D(
        mem_stage_inst_dmem_n4008), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__4_ ( .D(
        mem_stage_inst_dmem_n4009), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__5_ ( .D(
        mem_stage_inst_dmem_n4010), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__6_ ( .D(
        mem_stage_inst_dmem_n4011), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__7_ ( .D(
        mem_stage_inst_dmem_n4012), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__8_ ( .D(
        mem_stage_inst_dmem_n4013), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__9_ ( .D(
        mem_stage_inst_dmem_n4014), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__10_ ( .D(
        mem_stage_inst_dmem_n4015), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__11_ ( .D(
        mem_stage_inst_dmem_n4016), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__12_ ( .D(
        mem_stage_inst_dmem_n4017), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__13_ ( .D(
        mem_stage_inst_dmem_n4018), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__14_ ( .D(
        mem_stage_inst_dmem_n4019), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_215__15_ ( .D(
        mem_stage_inst_dmem_n4020), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_215__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__0_ ( .D(
        mem_stage_inst_dmem_n4069), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__1_ ( .D(
        mem_stage_inst_dmem_n4070), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__2_ ( .D(
        mem_stage_inst_dmem_n4071), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__3_ ( .D(
        mem_stage_inst_dmem_n4072), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__4_ ( .D(
        mem_stage_inst_dmem_n4073), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__5_ ( .D(
        mem_stage_inst_dmem_n4074), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__6_ ( .D(
        mem_stage_inst_dmem_n4075), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__7_ ( .D(
        mem_stage_inst_dmem_n4076), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__8_ ( .D(
        mem_stage_inst_dmem_n4077), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__9_ ( .D(
        mem_stage_inst_dmem_n4078), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__10_ ( .D(
        mem_stage_inst_dmem_n4079), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__11_ ( .D(
        mem_stage_inst_dmem_n4080), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__12_ ( .D(
        mem_stage_inst_dmem_n4081), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__13_ ( .D(
        mem_stage_inst_dmem_n4082), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__14_ ( .D(
        mem_stage_inst_dmem_n4083), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_219__15_ ( .D(
        mem_stage_inst_dmem_n4084), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_219__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__0_ ( .D(
        mem_stage_inst_dmem_n4133), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__1_ ( .D(
        mem_stage_inst_dmem_n4134), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__2_ ( .D(
        mem_stage_inst_dmem_n4135), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__3_ ( .D(
        mem_stage_inst_dmem_n4136), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__4_ ( .D(
        mem_stage_inst_dmem_n4137), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__5_ ( .D(
        mem_stage_inst_dmem_n4138), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__6_ ( .D(
        mem_stage_inst_dmem_n4139), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__7_ ( .D(
        mem_stage_inst_dmem_n4140), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__8_ ( .D(
        mem_stage_inst_dmem_n4141), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__9_ ( .D(
        mem_stage_inst_dmem_n4142), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__10_ ( .D(
        mem_stage_inst_dmem_n4143), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__11_ ( .D(
        mem_stage_inst_dmem_n4144), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__12_ ( .D(
        mem_stage_inst_dmem_n4145), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__13_ ( .D(
        mem_stage_inst_dmem_n4146), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__14_ ( .D(
        mem_stage_inst_dmem_n4147), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_223__15_ ( .D(
        mem_stage_inst_dmem_n4148), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_223__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__0_ ( .D(
        mem_stage_inst_dmem_n4197), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__1_ ( .D(
        mem_stage_inst_dmem_n4198), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__2_ ( .D(
        mem_stage_inst_dmem_n4199), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__3_ ( .D(
        mem_stage_inst_dmem_n4200), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__4_ ( .D(
        mem_stage_inst_dmem_n4201), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__5_ ( .D(
        mem_stage_inst_dmem_n4202), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__6_ ( .D(
        mem_stage_inst_dmem_n4203), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__7_ ( .D(
        mem_stage_inst_dmem_n4204), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__8_ ( .D(
        mem_stage_inst_dmem_n4205), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__9_ ( .D(
        mem_stage_inst_dmem_n4206), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__10_ ( .D(
        mem_stage_inst_dmem_n4207), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__11_ ( .D(
        mem_stage_inst_dmem_n4208), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__12_ ( .D(
        mem_stage_inst_dmem_n4209), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__13_ ( .D(
        mem_stage_inst_dmem_n4210), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__14_ ( .D(
        mem_stage_inst_dmem_n4211), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_227__15_ ( .D(
        mem_stage_inst_dmem_n4212), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_227__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__0_ ( .D(
        mem_stage_inst_dmem_n4261), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__1_ ( .D(
        mem_stage_inst_dmem_n4262), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__2_ ( .D(
        mem_stage_inst_dmem_n4263), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__3_ ( .D(
        mem_stage_inst_dmem_n4264), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__4_ ( .D(
        mem_stage_inst_dmem_n4265), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__5_ ( .D(
        mem_stage_inst_dmem_n4266), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__6_ ( .D(
        mem_stage_inst_dmem_n4267), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__7_ ( .D(
        mem_stage_inst_dmem_n4268), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__8_ ( .D(
        mem_stage_inst_dmem_n4269), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__9_ ( .D(
        mem_stage_inst_dmem_n4270), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__10_ ( .D(
        mem_stage_inst_dmem_n4271), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__11_ ( .D(
        mem_stage_inst_dmem_n4272), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__12_ ( .D(
        mem_stage_inst_dmem_n4273), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__13_ ( .D(
        mem_stage_inst_dmem_n4274), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__14_ ( .D(
        mem_stage_inst_dmem_n4275), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_231__15_ ( .D(
        mem_stage_inst_dmem_n4276), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_231__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__0_ ( .D(
        mem_stage_inst_dmem_n4325), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__1_ ( .D(
        mem_stage_inst_dmem_n4326), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__2_ ( .D(
        mem_stage_inst_dmem_n4327), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__3_ ( .D(
        mem_stage_inst_dmem_n4328), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__4_ ( .D(
        mem_stage_inst_dmem_n4329), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__5_ ( .D(
        mem_stage_inst_dmem_n4330), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__6_ ( .D(
        mem_stage_inst_dmem_n4331), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__7_ ( .D(
        mem_stage_inst_dmem_n4332), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__8_ ( .D(
        mem_stage_inst_dmem_n4333), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__9_ ( .D(
        mem_stage_inst_dmem_n4334), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__10_ ( .D(
        mem_stage_inst_dmem_n4335), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__11_ ( .D(
        mem_stage_inst_dmem_n4336), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__12_ ( .D(
        mem_stage_inst_dmem_n4337), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__13_ ( .D(
        mem_stage_inst_dmem_n4338), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__14_ ( .D(
        mem_stage_inst_dmem_n4339), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_235__15_ ( .D(
        mem_stage_inst_dmem_n4340), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_235__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__0_ ( .D(
        mem_stage_inst_dmem_n4389), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__1_ ( .D(
        mem_stage_inst_dmem_n4390), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__2_ ( .D(
        mem_stage_inst_dmem_n4391), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__3_ ( .D(
        mem_stage_inst_dmem_n4392), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__4_ ( .D(
        mem_stage_inst_dmem_n4393), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__5_ ( .D(
        mem_stage_inst_dmem_n4394), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__6_ ( .D(
        mem_stage_inst_dmem_n4395), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__7_ ( .D(
        mem_stage_inst_dmem_n4396), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__8_ ( .D(
        mem_stage_inst_dmem_n4397), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__9_ ( .D(
        mem_stage_inst_dmem_n4398), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__10_ ( .D(
        mem_stage_inst_dmem_n4399), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__11_ ( .D(
        mem_stage_inst_dmem_n4400), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__12_ ( .D(
        mem_stage_inst_dmem_n4401), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__13_ ( .D(
        mem_stage_inst_dmem_n4402), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__14_ ( .D(
        mem_stage_inst_dmem_n4403), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_239__15_ ( .D(
        mem_stage_inst_dmem_n4404), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_239__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__0_ ( .D(
        mem_stage_inst_dmem_n4453), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__1_ ( .D(
        mem_stage_inst_dmem_n4454), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__2_ ( .D(
        mem_stage_inst_dmem_n4455), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__3_ ( .D(
        mem_stage_inst_dmem_n4456), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__4_ ( .D(
        mem_stage_inst_dmem_n4457), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__5_ ( .D(
        mem_stage_inst_dmem_n4458), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__6_ ( .D(
        mem_stage_inst_dmem_n4459), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__7_ ( .D(
        mem_stage_inst_dmem_n4460), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__8_ ( .D(
        mem_stage_inst_dmem_n4461), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__9_ ( .D(
        mem_stage_inst_dmem_n4462), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__10_ ( .D(
        mem_stage_inst_dmem_n4463), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__11_ ( .D(
        mem_stage_inst_dmem_n4464), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__12_ ( .D(
        mem_stage_inst_dmem_n4465), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__13_ ( .D(
        mem_stage_inst_dmem_n4466), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__14_ ( .D(
        mem_stage_inst_dmem_n4467), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_243__15_ ( .D(
        mem_stage_inst_dmem_n4468), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_243__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__0_ ( .D(
        mem_stage_inst_dmem_n4517), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__1_ ( .D(
        mem_stage_inst_dmem_n4518), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__2_ ( .D(
        mem_stage_inst_dmem_n4519), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__3_ ( .D(
        mem_stage_inst_dmem_n4520), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__4_ ( .D(
        mem_stage_inst_dmem_n4521), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__5_ ( .D(
        mem_stage_inst_dmem_n4522), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__6_ ( .D(
        mem_stage_inst_dmem_n4523), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__7_ ( .D(
        mem_stage_inst_dmem_n4524), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__8_ ( .D(
        mem_stage_inst_dmem_n4525), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__9_ ( .D(
        mem_stage_inst_dmem_n4526), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__10_ ( .D(
        mem_stage_inst_dmem_n4527), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__11_ ( .D(
        mem_stage_inst_dmem_n4528), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__12_ ( .D(
        mem_stage_inst_dmem_n4529), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__13_ ( .D(
        mem_stage_inst_dmem_n4530), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__14_ ( .D(
        mem_stage_inst_dmem_n4531), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_247__15_ ( .D(
        mem_stage_inst_dmem_n4532), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_247__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__0_ ( .D(
        mem_stage_inst_dmem_n4581), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__1_ ( .D(
        mem_stage_inst_dmem_n4582), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__2_ ( .D(
        mem_stage_inst_dmem_n4583), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__3_ ( .D(
        mem_stage_inst_dmem_n4584), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__4_ ( .D(
        mem_stage_inst_dmem_n4585), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__5_ ( .D(
        mem_stage_inst_dmem_n4586), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__6_ ( .D(
        mem_stage_inst_dmem_n4587), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__7_ ( .D(
        mem_stage_inst_dmem_n4588), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__8_ ( .D(
        mem_stage_inst_dmem_n4589), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__9_ ( .D(
        mem_stage_inst_dmem_n4590), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__10_ ( .D(
        mem_stage_inst_dmem_n4591), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__11_ ( .D(
        mem_stage_inst_dmem_n4592), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__12_ ( .D(
        mem_stage_inst_dmem_n4593), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__13_ ( .D(
        mem_stage_inst_dmem_n4594), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__14_ ( .D(
        mem_stage_inst_dmem_n4595), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_251__15_ ( .D(
        mem_stage_inst_dmem_n4596), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_251__15_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__0_ ( .D(
        mem_stage_inst_dmem_n4645), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__0_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__1_ ( .D(
        mem_stage_inst_dmem_n4646), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__1_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__2_ ( .D(
        mem_stage_inst_dmem_n4647), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__2_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__3_ ( .D(
        mem_stage_inst_dmem_n4648), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__3_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__4_ ( .D(
        mem_stage_inst_dmem_n4649), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__4_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__5_ ( .D(
        mem_stage_inst_dmem_n4650), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__5_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__6_ ( .D(
        mem_stage_inst_dmem_n4651), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__6_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__7_ ( .D(
        mem_stage_inst_dmem_n4652), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__7_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__8_ ( .D(
        mem_stage_inst_dmem_n4653), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__8_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__9_ ( .D(
        mem_stage_inst_dmem_n4654), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__9_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__10_ ( .D(
        mem_stage_inst_dmem_n4655), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__10_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__11_ ( .D(
        mem_stage_inst_dmem_n4656), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__11_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__12_ ( .D(
        mem_stage_inst_dmem_n4657), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__12_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__13_ ( .D(
        mem_stage_inst_dmem_n4658), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__13_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__14_ ( .D(
        mem_stage_inst_dmem_n4659), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__14_) );
  DFFQ_X1M_A12TS mem_stage_inst_dmem_ram_reg_255__15_ ( .D(
        mem_stage_inst_dmem_n4660), .CK(clk), .Q(
        mem_stage_inst_dmem_ram_255__15_) );
  MXT2_X0P5M_A12TS wb_stage_inst_u16 ( .A(mem_pipeline_reg_out[21]), .B(
        mem_pipeline_reg_out[5]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[0]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u15 ( .A(mem_pipeline_reg_out[31]), .B(
        mem_pipeline_reg_out[15]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[10]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u14 ( .A(mem_pipeline_reg_out[32]), .B(
        mem_pipeline_reg_out[16]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[11]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u13 ( .A(mem_pipeline_reg_out[33]), .B(
        mem_pipeline_reg_out[17]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[12]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u12 ( .A(mem_pipeline_reg_out[34]), .B(
        mem_pipeline_reg_out[18]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[13]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u11 ( .A(mem_pipeline_reg_out[35]), .B(
        mem_pipeline_reg_out[19]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[14]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u10 ( .A(mem_pipeline_reg_out[36]), .B(
        mem_pipeline_reg_out[20]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[15]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u9 ( .A(mem_pipeline_reg_out[22]), .B(
        mem_pipeline_reg_out[6]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[1]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u8 ( .A(mem_pipeline_reg_out[23]), .B(
        mem_pipeline_reg_out[7]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[2]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u7 ( .A(mem_pipeline_reg_out[24]), .B(
        mem_pipeline_reg_out[8]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[3]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u6 ( .A(mem_pipeline_reg_out[25]), .B(
        mem_pipeline_reg_out[9]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[4]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u5 ( .A(mem_pipeline_reg_out[26]), .B(
        mem_pipeline_reg_out[10]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[5]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u4 ( .A(mem_pipeline_reg_out[27]), .B(
        mem_pipeline_reg_out[11]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[6]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u3 ( .A(mem_pipeline_reg_out[28]), .B(
        mem_pipeline_reg_out[12]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[7]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u2 ( .A(mem_pipeline_reg_out[29]), .B(
        mem_pipeline_reg_out[13]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[8]) );
  MXT2_X0P5M_A12TS wb_stage_inst_u1 ( .A(mem_pipeline_reg_out[30]), .B(
        mem_pipeline_reg_out[14]), .S0(mem_pipeline_reg_out[0]), .Y(
        reg_write_data[9]) );
  INV_X0P5B_A12TS register_file_inst_u271 ( .A(reg_write_dest[0]), .Y(
        register_file_inst_n199) );
  INV_X0P5B_A12TS register_file_inst_u270 ( .A(reg_write_dest[1]), .Y(
        register_file_inst_n201) );
  AND2_X0P5M_A12TS register_file_inst_u269 ( .A(reg_write_en), .B(
        reg_write_dest[2]), .Y(register_file_inst_n204) );
  AND3_X0P5M_A12TS register_file_inst_u268 ( .A(register_file_inst_n199), .B(
        register_file_inst_n201), .C(register_file_inst_n204), .Y(
        register_file_inst_n195) );
  MXT2_X0P5M_A12TS register_file_inst_u267 ( .A(
        register_file_inst_reg_array_4__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n100) );
  MXT2_X0P5M_A12TS register_file_inst_u266 ( .A(
        register_file_inst_reg_array_4__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n101) );
  MXT2_X0P5M_A12TS register_file_inst_u265 ( .A(
        register_file_inst_reg_array_4__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n102) );
  AND3_X0P5M_A12TS register_file_inst_u264 ( .A(register_file_inst_n204), .B(
        register_file_inst_n201), .C(reg_write_dest[0]), .Y(
        register_file_inst_n206) );
  MXT2_X0P5M_A12TS register_file_inst_u263 ( .A(
        register_file_inst_reg_array_5__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n103) );
  MXT2_X0P5M_A12TS register_file_inst_u262 ( .A(
        register_file_inst_reg_array_5__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n104) );
  MXT2_X0P5M_A12TS register_file_inst_u261 ( .A(
        register_file_inst_reg_array_5__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n105) );
  MXT2_X0P5M_A12TS register_file_inst_u260 ( .A(
        register_file_inst_reg_array_5__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n106) );
  MXT2_X0P5M_A12TS register_file_inst_u259 ( .A(
        register_file_inst_reg_array_5__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n107) );
  MXT2_X0P5M_A12TS register_file_inst_u258 ( .A(
        register_file_inst_reg_array_5__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n108) );
  MXT2_X0P5M_A12TS register_file_inst_u257 ( .A(
        register_file_inst_reg_array_5__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n109) );
  MXT2_X0P5M_A12TS register_file_inst_u256 ( .A(
        register_file_inst_reg_array_5__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n110) );
  MXT2_X0P5M_A12TS register_file_inst_u255 ( .A(
        register_file_inst_reg_array_5__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n111) );
  MXT2_X0P5M_A12TS register_file_inst_u254 ( .A(
        register_file_inst_reg_array_5__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n112) );
  MXT2_X0P5M_A12TS register_file_inst_u253 ( .A(
        register_file_inst_reg_array_5__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n113) );
  MXT2_X0P5M_A12TS register_file_inst_u252 ( .A(
        register_file_inst_reg_array_5__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n114) );
  MXT2_X0P5M_A12TS register_file_inst_u251 ( .A(
        register_file_inst_reg_array_5__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n115) );
  MXT2_X0P5M_A12TS register_file_inst_u250 ( .A(
        register_file_inst_reg_array_5__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n116) );
  MXT2_X0P5M_A12TS register_file_inst_u249 ( .A(
        register_file_inst_reg_array_5__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n117) );
  MXT2_X0P5M_A12TS register_file_inst_u248 ( .A(
        register_file_inst_reg_array_5__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n206), .Y(register_file_inst_n118) );
  AND3_X0P5M_A12TS register_file_inst_u247 ( .A(register_file_inst_n204), .B(
        register_file_inst_n199), .C(reg_write_dest[1]), .Y(
        register_file_inst_n205) );
  MXT2_X0P5M_A12TS register_file_inst_u246 ( .A(
        register_file_inst_reg_array_6__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n119) );
  MXT2_X0P5M_A12TS register_file_inst_u245 ( .A(
        register_file_inst_reg_array_6__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n120) );
  MXT2_X0P5M_A12TS register_file_inst_u244 ( .A(
        register_file_inst_reg_array_6__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n121) );
  MXT2_X0P5M_A12TS register_file_inst_u243 ( .A(
        register_file_inst_reg_array_6__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n122) );
  MXT2_X0P5M_A12TS register_file_inst_u242 ( .A(
        register_file_inst_reg_array_6__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n123) );
  MXT2_X0P5M_A12TS register_file_inst_u241 ( .A(
        register_file_inst_reg_array_6__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n124) );
  MXT2_X0P5M_A12TS register_file_inst_u240 ( .A(
        register_file_inst_reg_array_6__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n125) );
  MXT2_X0P5M_A12TS register_file_inst_u239 ( .A(
        register_file_inst_reg_array_6__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n126) );
  MXT2_X0P5M_A12TS register_file_inst_u238 ( .A(
        register_file_inst_reg_array_6__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n127) );
  MXT2_X0P5M_A12TS register_file_inst_u237 ( .A(
        register_file_inst_reg_array_6__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n128) );
  MXT2_X0P5M_A12TS register_file_inst_u236 ( .A(
        register_file_inst_reg_array_6__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n129) );
  MXT2_X0P5M_A12TS register_file_inst_u235 ( .A(
        register_file_inst_reg_array_6__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n130) );
  MXT2_X0P5M_A12TS register_file_inst_u234 ( .A(
        register_file_inst_reg_array_6__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n131) );
  MXT2_X0P5M_A12TS register_file_inst_u233 ( .A(
        register_file_inst_reg_array_6__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n132) );
  MXT2_X0P5M_A12TS register_file_inst_u232 ( .A(
        register_file_inst_reg_array_6__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n133) );
  MXT2_X0P5M_A12TS register_file_inst_u231 ( .A(
        register_file_inst_reg_array_6__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n205), .Y(register_file_inst_n134) );
  AND3_X0P5M_A12TS register_file_inst_u230 ( .A(reg_write_dest[0]), .B(
        register_file_inst_n204), .C(reg_write_dest[1]), .Y(
        register_file_inst_n203) );
  MXT2_X0P5M_A12TS register_file_inst_u229 ( .A(
        register_file_inst_reg_array_7__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n135) );
  MXT2_X0P5M_A12TS register_file_inst_u228 ( .A(
        register_file_inst_reg_array_7__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n136) );
  MXT2_X0P5M_A12TS register_file_inst_u227 ( .A(
        register_file_inst_reg_array_7__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n137) );
  MXT2_X0P5M_A12TS register_file_inst_u226 ( .A(
        register_file_inst_reg_array_7__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n138) );
  MXT2_X0P5M_A12TS register_file_inst_u225 ( .A(
        register_file_inst_reg_array_7__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n139) );
  MXT2_X0P5M_A12TS register_file_inst_u224 ( .A(
        register_file_inst_reg_array_7__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n140) );
  MXT2_X0P5M_A12TS register_file_inst_u223 ( .A(
        register_file_inst_reg_array_7__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n141) );
  MXT2_X0P5M_A12TS register_file_inst_u222 ( .A(
        register_file_inst_reg_array_7__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n142) );
  MXT2_X0P5M_A12TS register_file_inst_u221 ( .A(
        register_file_inst_reg_array_7__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n143) );
  MXT2_X0P5M_A12TS register_file_inst_u220 ( .A(
        register_file_inst_reg_array_7__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n144) );
  MXT2_X0P5M_A12TS register_file_inst_u219 ( .A(
        register_file_inst_reg_array_7__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n145) );
  MXT2_X0P5M_A12TS register_file_inst_u218 ( .A(
        register_file_inst_reg_array_7__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n146) );
  MXT2_X0P5M_A12TS register_file_inst_u217 ( .A(
        register_file_inst_reg_array_7__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n147) );
  MXT2_X0P5M_A12TS register_file_inst_u216 ( .A(
        register_file_inst_reg_array_7__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n148) );
  MXT2_X0P5M_A12TS register_file_inst_u215 ( .A(
        register_file_inst_reg_array_7__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n149) );
  MXT2_X0P5M_A12TS register_file_inst_u214 ( .A(
        register_file_inst_reg_array_7__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n203), .Y(register_file_inst_n150) );
  NOR2B_X0P5M_A12TS register_file_inst_u213 ( .AN(reg_write_en), .B(
        reg_write_dest[2]), .Y(register_file_inst_n197) );
  AND3_X0P5M_A12TS register_file_inst_u212 ( .A(register_file_inst_n199), .B(
        register_file_inst_n201), .C(register_file_inst_n197), .Y(
        register_file_inst_n202) );
  MXT2_X0P5M_A12TS register_file_inst_u211 ( .A(
        register_file_inst_reg_array_0__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n23) );
  MXT2_X0P5M_A12TS register_file_inst_u210 ( .A(
        register_file_inst_reg_array_0__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n24) );
  MXT2_X0P5M_A12TS register_file_inst_u209 ( .A(
        register_file_inst_reg_array_0__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n25) );
  MXT2_X0P5M_A12TS register_file_inst_u208 ( .A(
        register_file_inst_reg_array_0__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n26) );
  MXT2_X0P5M_A12TS register_file_inst_u207 ( .A(
        register_file_inst_reg_array_0__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n27) );
  MXT2_X0P5M_A12TS register_file_inst_u206 ( .A(
        register_file_inst_reg_array_0__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n28) );
  MXT2_X0P5M_A12TS register_file_inst_u205 ( .A(
        register_file_inst_reg_array_0__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n29) );
  MXT2_X0P5M_A12TS register_file_inst_u204 ( .A(
        register_file_inst_reg_array_0__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n30) );
  MXT2_X0P5M_A12TS register_file_inst_u203 ( .A(
        register_file_inst_reg_array_0__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n31) );
  MXT2_X0P5M_A12TS register_file_inst_u202 ( .A(
        register_file_inst_reg_array_0__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n32) );
  MXT2_X0P5M_A12TS register_file_inst_u201 ( .A(
        register_file_inst_reg_array_0__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n33) );
  MXT2_X0P5M_A12TS register_file_inst_u200 ( .A(
        register_file_inst_reg_array_0__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n34) );
  MXT2_X0P5M_A12TS register_file_inst_u199 ( .A(
        register_file_inst_reg_array_0__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n35) );
  MXT2_X0P5M_A12TS register_file_inst_u198 ( .A(
        register_file_inst_reg_array_0__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n36) );
  MXT2_X0P5M_A12TS register_file_inst_u197 ( .A(
        register_file_inst_reg_array_0__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n37) );
  MXT2_X0P5M_A12TS register_file_inst_u196 ( .A(
        register_file_inst_reg_array_0__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n202), .Y(register_file_inst_n38) );
  AND3_X0P5M_A12TS register_file_inst_u195 ( .A(register_file_inst_n197), .B(
        register_file_inst_n201), .C(reg_write_dest[0]), .Y(
        register_file_inst_n200) );
  MXT2_X0P5M_A12TS register_file_inst_u194 ( .A(
        register_file_inst_reg_array_1__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n39) );
  MXT2_X0P5M_A12TS register_file_inst_u193 ( .A(
        register_file_inst_reg_array_1__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n40) );
  MXT2_X0P5M_A12TS register_file_inst_u192 ( .A(
        register_file_inst_reg_array_1__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n41) );
  MXT2_X0P5M_A12TS register_file_inst_u191 ( .A(
        register_file_inst_reg_array_1__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n42) );
  MXT2_X0P5M_A12TS register_file_inst_u190 ( .A(
        register_file_inst_reg_array_1__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n43) );
  MXT2_X0P5M_A12TS register_file_inst_u189 ( .A(
        register_file_inst_reg_array_1__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n44) );
  MXT2_X0P5M_A12TS register_file_inst_u188 ( .A(
        register_file_inst_reg_array_1__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n45) );
  MXT2_X0P5M_A12TS register_file_inst_u187 ( .A(
        register_file_inst_reg_array_1__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n46) );
  MXT2_X0P5M_A12TS register_file_inst_u186 ( .A(
        register_file_inst_reg_array_1__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n47) );
  MXT2_X0P5M_A12TS register_file_inst_u185 ( .A(
        register_file_inst_reg_array_1__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n48) );
  MXT2_X0P5M_A12TS register_file_inst_u184 ( .A(
        register_file_inst_reg_array_1__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n49) );
  MXT2_X0P5M_A12TS register_file_inst_u183 ( .A(
        register_file_inst_reg_array_1__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n50) );
  MXT2_X0P5M_A12TS register_file_inst_u182 ( .A(
        register_file_inst_reg_array_1__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n51) );
  MXT2_X0P5M_A12TS register_file_inst_u181 ( .A(
        register_file_inst_reg_array_1__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n52) );
  MXT2_X0P5M_A12TS register_file_inst_u180 ( .A(
        register_file_inst_reg_array_1__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n53) );
  MXT2_X0P5M_A12TS register_file_inst_u179 ( .A(
        register_file_inst_reg_array_1__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n200), .Y(register_file_inst_n54) );
  AND3_X0P5M_A12TS register_file_inst_u178 ( .A(register_file_inst_n197), .B(
        register_file_inst_n199), .C(reg_write_dest[1]), .Y(
        register_file_inst_n198) );
  MXT2_X0P5M_A12TS register_file_inst_u177 ( .A(
        register_file_inst_reg_array_2__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n55) );
  MXT2_X0P5M_A12TS register_file_inst_u176 ( .A(
        register_file_inst_reg_array_2__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n56) );
  MXT2_X0P5M_A12TS register_file_inst_u175 ( .A(
        register_file_inst_reg_array_2__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n57) );
  MXT2_X0P5M_A12TS register_file_inst_u174 ( .A(
        register_file_inst_reg_array_2__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n58) );
  MXT2_X0P5M_A12TS register_file_inst_u173 ( .A(
        register_file_inst_reg_array_2__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n59) );
  MXT2_X0P5M_A12TS register_file_inst_u172 ( .A(
        register_file_inst_reg_array_2__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n60) );
  MXT2_X0P5M_A12TS register_file_inst_u171 ( .A(
        register_file_inst_reg_array_2__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n61) );
  MXT2_X0P5M_A12TS register_file_inst_u170 ( .A(
        register_file_inst_reg_array_2__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n62) );
  MXT2_X0P5M_A12TS register_file_inst_u169 ( .A(
        register_file_inst_reg_array_2__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n63) );
  MXT2_X0P5M_A12TS register_file_inst_u168 ( .A(
        register_file_inst_reg_array_2__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n64) );
  MXT2_X0P5M_A12TS register_file_inst_u167 ( .A(
        register_file_inst_reg_array_2__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n65) );
  MXT2_X0P5M_A12TS register_file_inst_u166 ( .A(
        register_file_inst_reg_array_2__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n66) );
  MXT2_X0P5M_A12TS register_file_inst_u165 ( .A(
        register_file_inst_reg_array_2__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n67) );
  MXT2_X0P5M_A12TS register_file_inst_u164 ( .A(
        register_file_inst_reg_array_2__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n68) );
  MXT2_X0P5M_A12TS register_file_inst_u163 ( .A(
        register_file_inst_reg_array_2__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n69) );
  MXT2_X0P5M_A12TS register_file_inst_u162 ( .A(
        register_file_inst_reg_array_2__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n198), .Y(register_file_inst_n70) );
  AND3_X0P5M_A12TS register_file_inst_u161 ( .A(reg_write_dest[0]), .B(
        register_file_inst_n197), .C(reg_write_dest[1]), .Y(
        register_file_inst_n196) );
  MXT2_X0P5M_A12TS register_file_inst_u160 ( .A(
        register_file_inst_reg_array_3__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n71) );
  MXT2_X0P5M_A12TS register_file_inst_u159 ( .A(
        register_file_inst_reg_array_3__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n72) );
  MXT2_X0P5M_A12TS register_file_inst_u158 ( .A(
        register_file_inst_reg_array_3__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n73) );
  MXT2_X0P5M_A12TS register_file_inst_u157 ( .A(
        register_file_inst_reg_array_3__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n74) );
  MXT2_X0P5M_A12TS register_file_inst_u156 ( .A(
        register_file_inst_reg_array_3__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n75) );
  MXT2_X0P5M_A12TS register_file_inst_u155 ( .A(
        register_file_inst_reg_array_3__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n76) );
  MXT2_X0P5M_A12TS register_file_inst_u154 ( .A(
        register_file_inst_reg_array_3__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n77) );
  MXT2_X0P5M_A12TS register_file_inst_u153 ( .A(
        register_file_inst_reg_array_3__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n78) );
  MXT2_X0P5M_A12TS register_file_inst_u152 ( .A(
        register_file_inst_reg_array_3__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n79) );
  MXT2_X0P5M_A12TS register_file_inst_u151 ( .A(
        register_file_inst_reg_array_3__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n80) );
  MXT2_X0P5M_A12TS register_file_inst_u150 ( .A(
        register_file_inst_reg_array_3__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n81) );
  MXT2_X0P5M_A12TS register_file_inst_u149 ( .A(
        register_file_inst_reg_array_3__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n82) );
  MXT2_X0P5M_A12TS register_file_inst_u148 ( .A(
        register_file_inst_reg_array_3__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n83) );
  MXT2_X0P5M_A12TS register_file_inst_u147 ( .A(
        register_file_inst_reg_array_3__13_), .B(reg_write_data[13]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n84) );
  MXT2_X0P5M_A12TS register_file_inst_u146 ( .A(
        register_file_inst_reg_array_3__14_), .B(reg_write_data[14]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n85) );
  MXT2_X0P5M_A12TS register_file_inst_u145 ( .A(
        register_file_inst_reg_array_3__15_), .B(reg_write_data[15]), .S0(
        register_file_inst_n196), .Y(register_file_inst_n86) );
  MXT2_X0P5M_A12TS register_file_inst_u144 ( .A(
        register_file_inst_reg_array_4__0_), .B(reg_write_data[0]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n87) );
  MXT2_X0P5M_A12TS register_file_inst_u143 ( .A(
        register_file_inst_reg_array_4__1_), .B(reg_write_data[1]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n88) );
  MXT2_X0P5M_A12TS register_file_inst_u142 ( .A(
        register_file_inst_reg_array_4__2_), .B(reg_write_data[2]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n89) );
  MXT2_X0P5M_A12TS register_file_inst_u141 ( .A(
        register_file_inst_reg_array_4__3_), .B(reg_write_data[3]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n90) );
  MXT2_X0P5M_A12TS register_file_inst_u140 ( .A(
        register_file_inst_reg_array_4__4_), .B(reg_write_data[4]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n91) );
  MXT2_X0P5M_A12TS register_file_inst_u139 ( .A(
        register_file_inst_reg_array_4__5_), .B(reg_write_data[5]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n92) );
  MXT2_X0P5M_A12TS register_file_inst_u138 ( .A(
        register_file_inst_reg_array_4__6_), .B(reg_write_data[6]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n93) );
  MXT2_X0P5M_A12TS register_file_inst_u137 ( .A(
        register_file_inst_reg_array_4__7_), .B(reg_write_data[7]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n94) );
  MXT2_X0P5M_A12TS register_file_inst_u136 ( .A(
        register_file_inst_reg_array_4__8_), .B(reg_write_data[8]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n95) );
  MXT2_X0P5M_A12TS register_file_inst_u135 ( .A(
        register_file_inst_reg_array_4__9_), .B(reg_write_data[9]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n96) );
  MXT2_X0P5M_A12TS register_file_inst_u134 ( .A(
        register_file_inst_reg_array_4__10_), .B(reg_write_data[10]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n97) );
  MXT2_X0P5M_A12TS register_file_inst_u133 ( .A(
        register_file_inst_reg_array_4__11_), .B(reg_write_data[11]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n98) );
  MXT2_X0P5M_A12TS register_file_inst_u132 ( .A(
        register_file_inst_reg_array_4__12_), .B(reg_write_data[12]), .S0(
        register_file_inst_n195), .Y(register_file_inst_n99) );
  OR3_X0P5M_A12TS register_file_inst_u131 ( .A(reg_read_addr_1[2]), .B(
        reg_read_addr_1[1]), .C(reg_read_addr_1[0]), .Y(
        register_file_inst_n194) );
  AND2_X0P5M_A12TS register_file_inst_u130 ( .A(register_file_inst_n440), .B(
        register_file_inst_n194), .Y(reg_read_data_1[0]) );
  AND2_X0P5M_A12TS register_file_inst_u129 ( .A(register_file_inst_n340), .B(
        register_file_inst_n194), .Y(reg_read_data_1[10]) );
  AND2_X0P5M_A12TS register_file_inst_u128 ( .A(register_file_inst_n330), .B(
        register_file_inst_n194), .Y(reg_read_data_1[11]) );
  AND2_X0P5M_A12TS register_file_inst_u127 ( .A(register_file_inst_n320), .B(
        register_file_inst_n194), .Y(reg_read_data_1[12]) );
  AND2_X0P5M_A12TS register_file_inst_u126 ( .A(register_file_inst_n310), .B(
        register_file_inst_n194), .Y(reg_read_data_1[13]) );
  AND2_X0P5M_A12TS register_file_inst_u125 ( .A(register_file_inst_n300), .B(
        register_file_inst_n194), .Y(reg_read_data_1[14]) );
  AND2_X0P5M_A12TS register_file_inst_u124 ( .A(register_file_inst_n290), .B(
        register_file_inst_n194), .Y(reg_read_data_1[15]) );
  AND2_X0P5M_A12TS register_file_inst_u123 ( .A(register_file_inst_n430), .B(
        register_file_inst_n194), .Y(reg_read_data_1[1]) );
  AND2_X0P5M_A12TS register_file_inst_u122 ( .A(register_file_inst_n420), .B(
        register_file_inst_n194), .Y(reg_read_data_1[2]) );
  AND2_X0P5M_A12TS register_file_inst_u121 ( .A(register_file_inst_n410), .B(
        register_file_inst_n194), .Y(reg_read_data_1[3]) );
  AND2_X0P5M_A12TS register_file_inst_u120 ( .A(register_file_inst_n400), .B(
        register_file_inst_n194), .Y(reg_read_data_1[4]) );
  AND2_X0P5M_A12TS register_file_inst_u119 ( .A(register_file_inst_n390), .B(
        register_file_inst_n194), .Y(reg_read_data_1[5]) );
  AND2_X0P5M_A12TS register_file_inst_u118 ( .A(register_file_inst_n380), .B(
        register_file_inst_n194), .Y(reg_read_data_1[6]) );
  AND2_X0P5M_A12TS register_file_inst_u117 ( .A(register_file_inst_n370), .B(
        register_file_inst_n194), .Y(reg_read_data_1[7]) );
  AND2_X0P5M_A12TS register_file_inst_u116 ( .A(register_file_inst_n360), .B(
        register_file_inst_n194), .Y(reg_read_data_1[8]) );
  AND2_X0P5M_A12TS register_file_inst_u115 ( .A(register_file_inst_n350), .B(
        register_file_inst_n194), .Y(reg_read_data_1[9]) );
  OR3_X0P5M_A12TS register_file_inst_u114 ( .A(reg_read_addr_2[2]), .B(
        reg_read_addr_2[1]), .C(reg_read_addr_2[0]), .Y(
        register_file_inst_n193) );
  AND2_X0P5M_A12TS register_file_inst_u113 ( .A(register_file_inst_n600), .B(
        register_file_inst_n193), .Y(reg_read_data_2[0]) );
  AND2_X0P5M_A12TS register_file_inst_u112 ( .A(register_file_inst_n500), .B(
        register_file_inst_n193), .Y(reg_read_data_2[10]) );
  AND2_X0P5M_A12TS register_file_inst_u111 ( .A(register_file_inst_n490), .B(
        register_file_inst_n193), .Y(reg_read_data_2[11]) );
  AND2_X0P5M_A12TS register_file_inst_u110 ( .A(register_file_inst_n480), .B(
        register_file_inst_n193), .Y(reg_read_data_2[12]) );
  AND2_X0P5M_A12TS register_file_inst_u109 ( .A(register_file_inst_n470), .B(
        register_file_inst_n193), .Y(reg_read_data_2[13]) );
  AND2_X0P5M_A12TS register_file_inst_u108 ( .A(register_file_inst_n460), .B(
        register_file_inst_n193), .Y(reg_read_data_2[14]) );
  AND2_X0P5M_A12TS register_file_inst_u107 ( .A(register_file_inst_n450), .B(
        register_file_inst_n193), .Y(reg_read_data_2[15]) );
  AND2_X0P5M_A12TS register_file_inst_u106 ( .A(register_file_inst_n590), .B(
        register_file_inst_n193), .Y(reg_read_data_2[1]) );
  AND2_X0P5M_A12TS register_file_inst_u105 ( .A(register_file_inst_n580), .B(
        register_file_inst_n193), .Y(reg_read_data_2[2]) );
  AND2_X0P5M_A12TS register_file_inst_u104 ( .A(register_file_inst_n570), .B(
        register_file_inst_n193), .Y(reg_read_data_2[3]) );
  AND2_X0P5M_A12TS register_file_inst_u103 ( .A(register_file_inst_n560), .B(
        register_file_inst_n193), .Y(reg_read_data_2[4]) );
  AND2_X0P5M_A12TS register_file_inst_u102 ( .A(register_file_inst_n550), .B(
        register_file_inst_n193), .Y(reg_read_data_2[5]) );
  AND2_X0P5M_A12TS register_file_inst_u101 ( .A(register_file_inst_n540), .B(
        register_file_inst_n193), .Y(reg_read_data_2[6]) );
  AND2_X0P5M_A12TS register_file_inst_u100 ( .A(register_file_inst_n530), .B(
        register_file_inst_n193), .Y(reg_read_data_2[7]) );
  AND2_X0P5M_A12TS register_file_inst_u99 ( .A(register_file_inst_n520), .B(
        register_file_inst_n193), .Y(reg_read_data_2[8]) );
  AND2_X0P5M_A12TS register_file_inst_u98 ( .A(register_file_inst_n510), .B(
        register_file_inst_n193), .Y(reg_read_data_2[9]) );
  MXT2_X1M_A12TS register_file_inst_u97 ( .A(register_file_inst_n165), .B(
        register_file_inst_n166), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n450) );
  MXT2_X1M_A12TS register_file_inst_u96 ( .A(register_file_inst_n163), .B(
        register_file_inst_n164), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n460) );
  MXT2_X1M_A12TS register_file_inst_u95 ( .A(register_file_inst_n161), .B(
        register_file_inst_n162), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n470) );
  MXT2_X1M_A12TS register_file_inst_u94 ( .A(register_file_inst_n159), .B(
        register_file_inst_n160), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n480) );
  MXT2_X1M_A12TS register_file_inst_u93 ( .A(register_file_inst_n157), .B(
        register_file_inst_n158), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n490) );
  MXT2_X1M_A12TS register_file_inst_u92 ( .A(register_file_inst_n155), .B(
        register_file_inst_n156), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n500) );
  MXT2_X1M_A12TS register_file_inst_u91 ( .A(register_file_inst_n153), .B(
        register_file_inst_n154), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n510) );
  MXT2_X1M_A12TS register_file_inst_u90 ( .A(register_file_inst_n151), .B(
        register_file_inst_n152), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n520) );
  MXT2_X1M_A12TS register_file_inst_u89 ( .A(register_file_inst_n21), .B(
        register_file_inst_n22), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n530) );
  MXT2_X1M_A12TS register_file_inst_u88 ( .A(register_file_inst_n19), .B(
        register_file_inst_n20), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n540) );
  MXIT4_X0P5M_A12TS register_file_inst_u87 ( .A(
        register_file_inst_reg_array_4__5_), .B(
        register_file_inst_reg_array_6__5_), .C(
        register_file_inst_reg_array_5__5_), .D(
        register_file_inst_reg_array_7__5_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n192) );
  MXIT4_X0P5M_A12TS register_file_inst_u86 ( .A(
        register_file_inst_reg_array_0__5_), .B(
        register_file_inst_reg_array_2__5_), .C(
        register_file_inst_reg_array_1__5_), .D(
        register_file_inst_reg_array_3__5_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n191) );
  MXIT2_X0P5M_A12TS register_file_inst_u85 ( .A(register_file_inst_n191), .B(
        register_file_inst_n192), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n550) );
  MXT4_X1M_A12TS register_file_inst_u84 ( .A(
        register_file_inst_reg_array_4__5_), .B(
        register_file_inst_reg_array_6__5_), .C(
        register_file_inst_reg_array_5__5_), .D(
        register_file_inst_reg_array_7__5_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n18) );
  MXT4_X1M_A12TS register_file_inst_u83 ( .A(
        register_file_inst_reg_array_0__5_), .B(
        register_file_inst_reg_array_2__5_), .C(
        register_file_inst_reg_array_1__5_), .D(
        register_file_inst_reg_array_3__5_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n17) );
  MXT2_X1M_A12TS register_file_inst_u82 ( .A(register_file_inst_n17), .B(
        register_file_inst_n18), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n390) );
  MXT4_X1M_A12TS register_file_inst_u81 ( .A(
        register_file_inst_reg_array_4__2_), .B(
        register_file_inst_reg_array_6__2_), .C(
        register_file_inst_reg_array_5__2_), .D(
        register_file_inst_reg_array_7__2_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n16) );
  MXT4_X1M_A12TS register_file_inst_u80 ( .A(
        register_file_inst_reg_array_0__2_), .B(
        register_file_inst_reg_array_2__2_), .C(
        register_file_inst_reg_array_1__2_), .D(
        register_file_inst_reg_array_3__2_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n15) );
  MXT2_X1M_A12TS register_file_inst_u79 ( .A(register_file_inst_n15), .B(
        register_file_inst_n16), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n420) );
  MXT4_X1M_A12TS register_file_inst_u78 ( .A(
        register_file_inst_reg_array_4__0_), .B(
        register_file_inst_reg_array_6__0_), .C(
        register_file_inst_reg_array_5__0_), .D(
        register_file_inst_reg_array_7__0_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n14) );
  MXT4_X1M_A12TS register_file_inst_u77 ( .A(
        register_file_inst_reg_array_0__0_), .B(
        register_file_inst_reg_array_2__0_), .C(
        register_file_inst_reg_array_1__0_), .D(
        register_file_inst_reg_array_3__0_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n13) );
  MXT2_X1M_A12TS register_file_inst_u76 ( .A(register_file_inst_n13), .B(
        register_file_inst_n14), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n440) );
  MXT4_X1M_A12TS register_file_inst_u75 ( .A(
        register_file_inst_reg_array_4__4_), .B(
        register_file_inst_reg_array_6__4_), .C(
        register_file_inst_reg_array_5__4_), .D(
        register_file_inst_reg_array_7__4_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n12) );
  MXT4_X1M_A12TS register_file_inst_u74 ( .A(
        register_file_inst_reg_array_0__4_), .B(
        register_file_inst_reg_array_2__4_), .C(
        register_file_inst_reg_array_1__4_), .D(
        register_file_inst_reg_array_3__4_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n11) );
  MXT2_X1M_A12TS register_file_inst_u73 ( .A(register_file_inst_n11), .B(
        register_file_inst_n12), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n400) );
  MXT4_X1M_A12TS register_file_inst_u72 ( .A(
        register_file_inst_reg_array_4__1_), .B(
        register_file_inst_reg_array_6__1_), .C(
        register_file_inst_reg_array_5__1_), .D(
        register_file_inst_reg_array_7__1_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n10) );
  MXT4_X1M_A12TS register_file_inst_u71 ( .A(
        register_file_inst_reg_array_0__1_), .B(
        register_file_inst_reg_array_2__1_), .C(
        register_file_inst_reg_array_1__1_), .D(
        register_file_inst_reg_array_3__1_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n9) );
  MXT2_X1M_A12TS register_file_inst_u70 ( .A(register_file_inst_n9), .B(
        register_file_inst_n10), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n430) );
  MXT4_X1M_A12TS register_file_inst_u69 ( .A(
        register_file_inst_reg_array_4__14_), .B(
        register_file_inst_reg_array_6__14_), .C(
        register_file_inst_reg_array_5__14_), .D(
        register_file_inst_reg_array_7__14_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n8) );
  MXT4_X1M_A12TS register_file_inst_u68 ( .A(
        register_file_inst_reg_array_0__14_), .B(
        register_file_inst_reg_array_2__14_), .C(
        register_file_inst_reg_array_1__14_), .D(
        register_file_inst_reg_array_3__14_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n7) );
  MXT2_X1M_A12TS register_file_inst_u67 ( .A(register_file_inst_n7), .B(
        register_file_inst_n8), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n300) );
  MXT4_X1M_A12TS register_file_inst_u66 ( .A(
        register_file_inst_reg_array_4__12_), .B(
        register_file_inst_reg_array_6__12_), .C(
        register_file_inst_reg_array_5__12_), .D(
        register_file_inst_reg_array_7__12_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n6) );
  MXT4_X1M_A12TS register_file_inst_u65 ( .A(
        register_file_inst_reg_array_0__12_), .B(
        register_file_inst_reg_array_2__12_), .C(
        register_file_inst_reg_array_1__12_), .D(
        register_file_inst_reg_array_3__12_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n5) );
  MXT2_X1M_A12TS register_file_inst_u64 ( .A(register_file_inst_n5), .B(
        register_file_inst_n6), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n320) );
  MXT4_X1M_A12TS register_file_inst_u63 ( .A(
        register_file_inst_reg_array_4__8_), .B(
        register_file_inst_reg_array_6__8_), .C(
        register_file_inst_reg_array_5__8_), .D(
        register_file_inst_reg_array_7__8_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n4) );
  MXT4_X1M_A12TS register_file_inst_u62 ( .A(
        register_file_inst_reg_array_0__8_), .B(
        register_file_inst_reg_array_2__8_), .C(
        register_file_inst_reg_array_1__8_), .D(
        register_file_inst_reg_array_3__8_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n3) );
  MXT2_X1M_A12TS register_file_inst_u61 ( .A(register_file_inst_n3), .B(
        register_file_inst_n4), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n360) );
  MXIT4_X0P7M_A12TS register_file_inst_u60 ( .A(
        register_file_inst_reg_array_4__15_), .B(
        register_file_inst_reg_array_6__15_), .C(
        register_file_inst_reg_array_5__15_), .D(
        register_file_inst_reg_array_7__15_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n180) );
  MXIT4_X0P7M_A12TS register_file_inst_u59 ( .A(
        register_file_inst_reg_array_0__15_), .B(
        register_file_inst_reg_array_2__15_), .C(
        register_file_inst_reg_array_1__15_), .D(
        register_file_inst_reg_array_3__15_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n179) );
  MXIT2_X0P7M_A12TS register_file_inst_u58 ( .A(register_file_inst_n179), .B(
        register_file_inst_n180), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n290) );
  MXIT4_X0P7M_A12TS register_file_inst_u57 ( .A(
        register_file_inst_reg_array_4__13_), .B(
        register_file_inst_reg_array_6__13_), .C(
        register_file_inst_reg_array_5__13_), .D(
        register_file_inst_reg_array_7__13_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n178) );
  MXIT4_X0P7M_A12TS register_file_inst_u56 ( .A(
        register_file_inst_reg_array_0__13_), .B(
        register_file_inst_reg_array_2__13_), .C(
        register_file_inst_reg_array_1__13_), .D(
        register_file_inst_reg_array_3__13_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n177) );
  MXIT2_X0P7M_A12TS register_file_inst_u55 ( .A(register_file_inst_n177), .B(
        register_file_inst_n178), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n310) );
  MXT4_X1M_A12TS register_file_inst_u54 ( .A(
        register_file_inst_reg_array_4__9_), .B(
        register_file_inst_reg_array_6__9_), .C(
        register_file_inst_reg_array_5__9_), .D(
        register_file_inst_reg_array_7__9_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n2) );
  MXT4_X1M_A12TS register_file_inst_u53 ( .A(
        register_file_inst_reg_array_0__9_), .B(
        register_file_inst_reg_array_2__9_), .C(
        register_file_inst_reg_array_1__9_), .D(
        register_file_inst_reg_array_3__9_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n1) );
  MXT2_X1M_A12TS register_file_inst_u52 ( .A(register_file_inst_n1), .B(
        register_file_inst_n2), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n350) );
  MXIT4_X0P7M_A12TS register_file_inst_u51 ( .A(
        register_file_inst_reg_array_4__10_), .B(
        register_file_inst_reg_array_6__10_), .C(
        register_file_inst_reg_array_5__10_), .D(
        register_file_inst_reg_array_7__10_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n174) );
  MXIT4_X0P7M_A12TS register_file_inst_u50 ( .A(
        register_file_inst_reg_array_0__10_), .B(
        register_file_inst_reg_array_2__10_), .C(
        register_file_inst_reg_array_1__10_), .D(
        register_file_inst_reg_array_3__10_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n173) );
  MXIT2_X0P7M_A12TS register_file_inst_u49 ( .A(register_file_inst_n173), .B(
        register_file_inst_n174), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n340) );
  MXIT4_X0P7M_A12TS register_file_inst_u48 ( .A(
        register_file_inst_reg_array_4__6_), .B(
        register_file_inst_reg_array_6__6_), .C(
        register_file_inst_reg_array_5__6_), .D(
        register_file_inst_reg_array_7__6_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n170) );
  MXIT4_X0P7M_A12TS register_file_inst_u47 ( .A(
        register_file_inst_reg_array_0__6_), .B(
        register_file_inst_reg_array_2__6_), .C(
        register_file_inst_reg_array_1__6_), .D(
        register_file_inst_reg_array_3__6_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n169) );
  MXIT2_X0P7M_A12TS register_file_inst_u46 ( .A(register_file_inst_n169), .B(
        register_file_inst_n170), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n380) );
  MXIT4_X0P7M_A12TS register_file_inst_u45 ( .A(
        register_file_inst_reg_array_4__3_), .B(
        register_file_inst_reg_array_6__3_), .C(
        register_file_inst_reg_array_5__3_), .D(
        register_file_inst_reg_array_7__3_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n168) );
  MXIT4_X0P7M_A12TS register_file_inst_u44 ( .A(
        register_file_inst_reg_array_0__3_), .B(
        register_file_inst_reg_array_2__3_), .C(
        register_file_inst_reg_array_1__3_), .D(
        register_file_inst_reg_array_3__3_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n167) );
  MXIT2_X0P7M_A12TS register_file_inst_u43 ( .A(register_file_inst_n167), .B(
        register_file_inst_n168), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n410) );
  MXIT4_X0P5M_A12TS register_file_inst_u42 ( .A(
        register_file_inst_reg_array_4__4_), .B(
        register_file_inst_reg_array_6__4_), .C(
        register_file_inst_reg_array_5__4_), .D(
        register_file_inst_reg_array_7__4_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n190) );
  MXIT4_X0P5M_A12TS register_file_inst_u41 ( .A(
        register_file_inst_reg_array_0__4_), .B(
        register_file_inst_reg_array_2__4_), .C(
        register_file_inst_reg_array_1__4_), .D(
        register_file_inst_reg_array_3__4_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n189) );
  MXIT2_X0P5M_A12TS register_file_inst_u40 ( .A(register_file_inst_n189), .B(
        register_file_inst_n190), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n560) );
  MXIT4_X0P5M_A12TS register_file_inst_u39 ( .A(
        register_file_inst_reg_array_4__3_), .B(
        register_file_inst_reg_array_6__3_), .C(
        register_file_inst_reg_array_5__3_), .D(
        register_file_inst_reg_array_7__3_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n188) );
  MXIT4_X0P5M_A12TS register_file_inst_u38 ( .A(
        register_file_inst_reg_array_0__3_), .B(
        register_file_inst_reg_array_2__3_), .C(
        register_file_inst_reg_array_1__3_), .D(
        register_file_inst_reg_array_3__3_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n187) );
  MXIT2_X0P7M_A12TS register_file_inst_u37 ( .A(register_file_inst_n187), .B(
        register_file_inst_n188), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n570) );
  MXIT4_X0P5M_A12TS register_file_inst_u36 ( .A(
        register_file_inst_reg_array_4__2_), .B(
        register_file_inst_reg_array_6__2_), .C(
        register_file_inst_reg_array_5__2_), .D(
        register_file_inst_reg_array_7__2_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n186) );
  MXIT4_X0P5M_A12TS register_file_inst_u35 ( .A(
        register_file_inst_reg_array_0__2_), .B(
        register_file_inst_reg_array_2__2_), .C(
        register_file_inst_reg_array_1__2_), .D(
        register_file_inst_reg_array_3__2_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n185) );
  MXIT2_X0P7M_A12TS register_file_inst_u34 ( .A(register_file_inst_n185), .B(
        register_file_inst_n186), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n580) );
  MXIT4_X0P5M_A12TS register_file_inst_u33 ( .A(
        register_file_inst_reg_array_4__1_), .B(
        register_file_inst_reg_array_6__1_), .C(
        register_file_inst_reg_array_5__1_), .D(
        register_file_inst_reg_array_7__1_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n184) );
  MXIT4_X0P5M_A12TS register_file_inst_u32 ( .A(
        register_file_inst_reg_array_0__1_), .B(
        register_file_inst_reg_array_2__1_), .C(
        register_file_inst_reg_array_1__1_), .D(
        register_file_inst_reg_array_3__1_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n183) );
  MXIT2_X0P7M_A12TS register_file_inst_u31 ( .A(register_file_inst_n183), .B(
        register_file_inst_n184), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n590) );
  MXIT4_X0P5M_A12TS register_file_inst_u30 ( .A(
        register_file_inst_reg_array_4__0_), .B(
        register_file_inst_reg_array_6__0_), .C(
        register_file_inst_reg_array_5__0_), .D(
        register_file_inst_reg_array_7__0_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n182) );
  MXIT4_X0P5M_A12TS register_file_inst_u29 ( .A(
        register_file_inst_reg_array_0__0_), .B(
        register_file_inst_reg_array_2__0_), .C(
        register_file_inst_reg_array_1__0_), .D(
        register_file_inst_reg_array_3__0_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n181) );
  MXIT2_X0P7M_A12TS register_file_inst_u28 ( .A(register_file_inst_n181), .B(
        register_file_inst_n182), .S0(reg_read_addr_2[2]), .Y(
        register_file_inst_n600) );
  MXIT4_X0P7M_A12TS register_file_inst_u27 ( .A(
        register_file_inst_reg_array_4__11_), .B(
        register_file_inst_reg_array_6__11_), .C(
        register_file_inst_reg_array_5__11_), .D(
        register_file_inst_reg_array_7__11_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n176) );
  MXIT4_X0P7M_A12TS register_file_inst_u26 ( .A(
        register_file_inst_reg_array_0__11_), .B(
        register_file_inst_reg_array_2__11_), .C(
        register_file_inst_reg_array_1__11_), .D(
        register_file_inst_reg_array_3__11_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n175) );
  MXIT2_X0P7M_A12TS register_file_inst_u25 ( .A(register_file_inst_n175), .B(
        register_file_inst_n176), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n330) );
  MXIT4_X0P7M_A12TS register_file_inst_u24 ( .A(
        register_file_inst_reg_array_4__7_), .B(
        register_file_inst_reg_array_6__7_), .C(
        register_file_inst_reg_array_5__7_), .D(
        register_file_inst_reg_array_7__7_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n172) );
  MXIT4_X0P7M_A12TS register_file_inst_u23 ( .A(
        register_file_inst_reg_array_0__7_), .B(
        register_file_inst_reg_array_2__7_), .C(
        register_file_inst_reg_array_1__7_), .D(
        register_file_inst_reg_array_3__7_), .S0(reg_read_addr_1[1]), .S1(
        reg_read_addr_1[0]), .Y(register_file_inst_n171) );
  MXIT2_X0P7M_A12TS register_file_inst_u22 ( .A(register_file_inst_n171), .B(
        register_file_inst_n172), .S0(reg_read_addr_1[2]), .Y(
        register_file_inst_n370) );
  MXT4_X0P5M_A12TS register_file_inst_u21 ( .A(
        register_file_inst_reg_array_0__15_), .B(
        register_file_inst_reg_array_2__15_), .C(
        register_file_inst_reg_array_1__15_), .D(
        register_file_inst_reg_array_3__15_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n165) );
  MXT4_X0P5M_A12TS register_file_inst_u20 ( .A(
        register_file_inst_reg_array_4__15_), .B(
        register_file_inst_reg_array_6__15_), .C(
        register_file_inst_reg_array_5__15_), .D(
        register_file_inst_reg_array_7__15_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n166) );
  MXT4_X0P5M_A12TS register_file_inst_u19 ( .A(
        register_file_inst_reg_array_0__14_), .B(
        register_file_inst_reg_array_2__14_), .C(
        register_file_inst_reg_array_1__14_), .D(
        register_file_inst_reg_array_3__14_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n163) );
  MXT4_X0P5M_A12TS register_file_inst_u18 ( .A(
        register_file_inst_reg_array_4__14_), .B(
        register_file_inst_reg_array_6__14_), .C(
        register_file_inst_reg_array_5__14_), .D(
        register_file_inst_reg_array_7__14_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n164) );
  MXT4_X0P5M_A12TS register_file_inst_u17 ( .A(
        register_file_inst_reg_array_0__13_), .B(
        register_file_inst_reg_array_2__13_), .C(
        register_file_inst_reg_array_1__13_), .D(
        register_file_inst_reg_array_3__13_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n161) );
  MXT4_X0P5M_A12TS register_file_inst_u16 ( .A(
        register_file_inst_reg_array_4__13_), .B(
        register_file_inst_reg_array_6__13_), .C(
        register_file_inst_reg_array_5__13_), .D(
        register_file_inst_reg_array_7__13_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n162) );
  MXT4_X0P5M_A12TS register_file_inst_u15 ( .A(
        register_file_inst_reg_array_0__12_), .B(
        register_file_inst_reg_array_2__12_), .C(
        register_file_inst_reg_array_1__12_), .D(
        register_file_inst_reg_array_3__12_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n159) );
  MXT4_X0P5M_A12TS register_file_inst_u14 ( .A(
        register_file_inst_reg_array_4__12_), .B(
        register_file_inst_reg_array_6__12_), .C(
        register_file_inst_reg_array_5__12_), .D(
        register_file_inst_reg_array_7__12_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n160) );
  MXT4_X0P5M_A12TS register_file_inst_u13 ( .A(
        register_file_inst_reg_array_0__11_), .B(
        register_file_inst_reg_array_2__11_), .C(
        register_file_inst_reg_array_1__11_), .D(
        register_file_inst_reg_array_3__11_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n157) );
  MXT4_X0P5M_A12TS register_file_inst_u12 ( .A(
        register_file_inst_reg_array_4__11_), .B(
        register_file_inst_reg_array_6__11_), .C(
        register_file_inst_reg_array_5__11_), .D(
        register_file_inst_reg_array_7__11_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n158) );
  MXT4_X0P5M_A12TS register_file_inst_u11 ( .A(
        register_file_inst_reg_array_0__10_), .B(
        register_file_inst_reg_array_2__10_), .C(
        register_file_inst_reg_array_1__10_), .D(
        register_file_inst_reg_array_3__10_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n155) );
  MXT4_X0P5M_A12TS register_file_inst_u10 ( .A(
        register_file_inst_reg_array_4__10_), .B(
        register_file_inst_reg_array_6__10_), .C(
        register_file_inst_reg_array_5__10_), .D(
        register_file_inst_reg_array_7__10_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n156) );
  MXT4_X0P5M_A12TS register_file_inst_u9 ( .A(
        register_file_inst_reg_array_0__9_), .B(
        register_file_inst_reg_array_2__9_), .C(
        register_file_inst_reg_array_1__9_), .D(
        register_file_inst_reg_array_3__9_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n153) );
  MXT4_X0P5M_A12TS register_file_inst_u8 ( .A(
        register_file_inst_reg_array_4__9_), .B(
        register_file_inst_reg_array_6__9_), .C(
        register_file_inst_reg_array_5__9_), .D(
        register_file_inst_reg_array_7__9_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n154) );
  MXT4_X0P5M_A12TS register_file_inst_u7 ( .A(
        register_file_inst_reg_array_0__8_), .B(
        register_file_inst_reg_array_2__8_), .C(
        register_file_inst_reg_array_1__8_), .D(
        register_file_inst_reg_array_3__8_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n151) );
  MXT4_X0P5M_A12TS register_file_inst_u6 ( .A(
        register_file_inst_reg_array_4__8_), .B(
        register_file_inst_reg_array_6__8_), .C(
        register_file_inst_reg_array_5__8_), .D(
        register_file_inst_reg_array_7__8_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n152) );
  MXT4_X0P5M_A12TS register_file_inst_u5 ( .A(
        register_file_inst_reg_array_0__7_), .B(
        register_file_inst_reg_array_2__7_), .C(
        register_file_inst_reg_array_1__7_), .D(
        register_file_inst_reg_array_3__7_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n21) );
  MXT4_X0P5M_A12TS register_file_inst_u4 ( .A(
        register_file_inst_reg_array_4__7_), .B(
        register_file_inst_reg_array_6__7_), .C(
        register_file_inst_reg_array_5__7_), .D(
        register_file_inst_reg_array_7__7_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n22) );
  MXT4_X0P5M_A12TS register_file_inst_u3 ( .A(
        register_file_inst_reg_array_0__6_), .B(
        register_file_inst_reg_array_2__6_), .C(
        register_file_inst_reg_array_1__6_), .D(
        register_file_inst_reg_array_3__6_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n19) );
  MXT4_X0P5M_A12TS register_file_inst_u2 ( .A(
        register_file_inst_reg_array_4__6_), .B(
        register_file_inst_reg_array_6__6_), .C(
        register_file_inst_reg_array_5__6_), .D(
        register_file_inst_reg_array_7__6_), .S0(reg_read_addr_2[1]), .S1(
        reg_read_addr_2[0]), .Y(register_file_inst_n20) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__0_ ( .D(
        register_file_inst_n55), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__1_ ( .D(
        register_file_inst_n56), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__2_ ( .D(
        register_file_inst_n57), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__3_ ( .D(
        register_file_inst_n58), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__4_ ( .D(
        register_file_inst_n59), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__5_ ( .D(
        register_file_inst_n60), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__6_ ( .D(
        register_file_inst_n61), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__7_ ( .D(
        register_file_inst_n62), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__8_ ( .D(
        register_file_inst_n63), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__9_ ( .D(
        register_file_inst_n64), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__10_ ( .D(
        register_file_inst_n65), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__11_ ( .D(
        register_file_inst_n66), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__12_ ( .D(
        register_file_inst_n67), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__13_ ( .D(
        register_file_inst_n68), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__14_ ( .D(
        register_file_inst_n69), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_2__15_ ( .D(
        register_file_inst_n70), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_2__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__0_ ( .D(
        register_file_inst_n119), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__1_ ( .D(
        register_file_inst_n120), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__2_ ( .D(
        register_file_inst_n121), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__3_ ( .D(
        register_file_inst_n122), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__4_ ( .D(
        register_file_inst_n123), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__5_ ( .D(
        register_file_inst_n124), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__6_ ( .D(
        register_file_inst_n125), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__7_ ( .D(
        register_file_inst_n126), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__8_ ( .D(
        register_file_inst_n127), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__9_ ( .D(
        register_file_inst_n128), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__10_ ( .D(
        register_file_inst_n129), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__11_ ( .D(
        register_file_inst_n130), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__12_ ( .D(
        register_file_inst_n131), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__13_ ( .D(
        register_file_inst_n132), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__14_ ( .D(
        register_file_inst_n133), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_6__15_ ( .D(
        register_file_inst_n134), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_6__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__0_ ( .D(
        register_file_inst_n23), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__1_ ( .D(
        register_file_inst_n24), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__2_ ( .D(
        register_file_inst_n25), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__3_ ( .D(
        register_file_inst_n26), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__4_ ( .D(
        register_file_inst_n27), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__5_ ( .D(
        register_file_inst_n28), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__6_ ( .D(
        register_file_inst_n29), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__7_ ( .D(
        register_file_inst_n30), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__8_ ( .D(
        register_file_inst_n31), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__9_ ( .D(
        register_file_inst_n32), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__10_ ( .D(
        register_file_inst_n33), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__11_ ( .D(
        register_file_inst_n34), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__12_ ( .D(
        register_file_inst_n35), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__13_ ( .D(
        register_file_inst_n36), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__14_ ( .D(
        register_file_inst_n37), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_0__15_ ( .D(
        register_file_inst_n38), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_0__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__0_ ( .D(
        register_file_inst_n87), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__1_ ( .D(
        register_file_inst_n88), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__2_ ( .D(
        register_file_inst_n89), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__3_ ( .D(
        register_file_inst_n90), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__4_ ( .D(
        register_file_inst_n91), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__5_ ( .D(
        register_file_inst_n92), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__6_ ( .D(
        register_file_inst_n93), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__7_ ( .D(
        register_file_inst_n94), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__8_ ( .D(
        register_file_inst_n95), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__9_ ( .D(
        register_file_inst_n96), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__10_ ( .D(
        register_file_inst_n97), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__11_ ( .D(
        register_file_inst_n98), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__12_ ( .D(
        register_file_inst_n99), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__13_ ( .D(
        register_file_inst_n100), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__14_ ( .D(
        register_file_inst_n101), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_4__15_ ( .D(
        register_file_inst_n102), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_4__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__0_ ( .D(
        register_file_inst_n39), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__1_ ( .D(
        register_file_inst_n40), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__2_ ( .D(
        register_file_inst_n41), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__3_ ( .D(
        register_file_inst_n42), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__4_ ( .D(
        register_file_inst_n43), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__5_ ( .D(
        register_file_inst_n44), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__6_ ( .D(
        register_file_inst_n45), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__7_ ( .D(
        register_file_inst_n46), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__8_ ( .D(
        register_file_inst_n47), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__9_ ( .D(
        register_file_inst_n48), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__10_ ( .D(
        register_file_inst_n49), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__11_ ( .D(
        register_file_inst_n50), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__12_ ( .D(
        register_file_inst_n51), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__13_ ( .D(
        register_file_inst_n52), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__14_ ( .D(
        register_file_inst_n53), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_1__15_ ( .D(
        register_file_inst_n54), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_1__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__0_ ( .D(
        register_file_inst_n103), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__1_ ( .D(
        register_file_inst_n104), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__2_ ( .D(
        register_file_inst_n105), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__3_ ( .D(
        register_file_inst_n106), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__4_ ( .D(
        register_file_inst_n107), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__5_ ( .D(
        register_file_inst_n108), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__6_ ( .D(
        register_file_inst_n109), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__7_ ( .D(
        register_file_inst_n110), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__8_ ( .D(
        register_file_inst_n111), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__9_ ( .D(
        register_file_inst_n112), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__10_ ( .D(
        register_file_inst_n113), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__11_ ( .D(
        register_file_inst_n114), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__12_ ( .D(
        register_file_inst_n115), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__13_ ( .D(
        register_file_inst_n116), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__14_ ( .D(
        register_file_inst_n117), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_5__15_ ( .D(
        register_file_inst_n118), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_5__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__0_ ( .D(
        register_file_inst_n71), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__1_ ( .D(
        register_file_inst_n72), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__2_ ( .D(
        register_file_inst_n73), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__3_ ( .D(
        register_file_inst_n74), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__4_ ( .D(
        register_file_inst_n75), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__5_ ( .D(
        register_file_inst_n76), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__6_ ( .D(
        register_file_inst_n77), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__7_ ( .D(
        register_file_inst_n78), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__8_ ( .D(
        register_file_inst_n79), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__9_ ( .D(
        register_file_inst_n80), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__10_ ( .D(
        register_file_inst_n81), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__11_ ( .D(
        register_file_inst_n82), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__12_ ( .D(
        register_file_inst_n83), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__13_ ( .D(
        register_file_inst_n84), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__14_ ( .D(
        register_file_inst_n85), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_3__15_ ( .D(
        register_file_inst_n86), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_3__15_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__0_ ( .D(
        register_file_inst_n135), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__0_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__1_ ( .D(
        register_file_inst_n136), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__1_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__2_ ( .D(
        register_file_inst_n137), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__2_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__3_ ( .D(
        register_file_inst_n138), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__3_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__4_ ( .D(
        register_file_inst_n139), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__4_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__5_ ( .D(
        register_file_inst_n140), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__5_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__6_ ( .D(
        register_file_inst_n141), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__6_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__7_ ( .D(
        register_file_inst_n142), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__7_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__8_ ( .D(
        register_file_inst_n143), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__8_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__9_ ( .D(
        register_file_inst_n144), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__9_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__10_ ( .D(
        register_file_inst_n145), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__10_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__11_ ( .D(
        register_file_inst_n146), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__11_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__12_ ( .D(
        register_file_inst_n147), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__12_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__13_ ( .D(
        register_file_inst_n148), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__13_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__14_ ( .D(
        register_file_inst_n149), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__14_) );
  DFFRPQ_X1M_A12TS register_file_inst_reg_array_reg_7__15_ ( .D(
        register_file_inst_n150), .CK(clk), .R(rst), .Q(
        register_file_inst_reg_array_7__15_) );
  INV_X0P5B_A12TS hazard_detection_unit_inst_u34 ( .A(reg_read_addr_1[1]), .Y(
        hazard_detection_unit_inst_n18) );
  INV_X0P5B_A12TS hazard_detection_unit_inst_u33 ( .A(reg_read_addr_1[2]), .Y(
        hazard_detection_unit_inst_n19) );
  INV_X0P5B_A12TS hazard_detection_unit_inst_u32 ( .A(reg_read_addr_1[0]), .Y(
        hazard_detection_unit_inst_n20) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u31 ( .A(mem_op_dest[0]), .B(
        reg_read_addr_1[0]), .Y(hazard_detection_unit_inst_n26) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u30 ( .A(mem_op_dest[2]), .B(
        reg_read_addr_1[2]), .Y(hazard_detection_unit_inst_n27) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u29 ( .A(mem_op_dest[1]), .B(
        reg_read_addr_1[1]), .Y(hazard_detection_unit_inst_n28) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u28 ( .A(ex_op_dest[2]), .B(
        hazard_detection_unit_inst_n19), .Y(hazard_detection_unit_inst_n31) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u27 ( .A(ex_op_dest[0]), .B(
        hazard_detection_unit_inst_n20), .Y(hazard_detection_unit_inst_n32) );
  NOR2_X0P5A_A12TS hazard_detection_unit_inst_u26 ( .A(
        hazard_detection_unit_inst_n31), .B(hazard_detection_unit_inst_n32), 
        .Y(hazard_detection_unit_inst_n29) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u25 ( .A(ex_op_dest[1]), .B(
        reg_read_addr_1[1]), .Y(hazard_detection_unit_inst_n30) );
  AOI32_X0P5M_A12TS hazard_detection_unit_inst_u24 ( .A0(
        hazard_detection_unit_inst_n26), .A1(hazard_detection_unit_inst_n27), 
        .A2(hazard_detection_unit_inst_n28), .B0(
        hazard_detection_unit_inst_n29), .B1(hazard_detection_unit_inst_n30), 
        .Y(hazard_detection_unit_inst_n21) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u23 ( .A(reg_write_dest[0]), 
        .B(reg_read_addr_1[0]), .Y(hazard_detection_unit_inst_n23) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u22 ( .A(reg_write_dest[2]), 
        .B(reg_read_addr_1[2]), .Y(hazard_detection_unit_inst_n24) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u21 ( .A(reg_write_dest[1]), 
        .B(reg_read_addr_1[1]), .Y(hazard_detection_unit_inst_n25) );
  NAND3_X0P5A_A12TS hazard_detection_unit_inst_u20 ( .A(
        hazard_detection_unit_inst_n23), .B(hazard_detection_unit_inst_n24), 
        .C(hazard_detection_unit_inst_n25), .Y(hazard_detection_unit_inst_n22)
         );
  AOI32_X0P5M_A12TS hazard_detection_unit_inst_u19 ( .A0(
        hazard_detection_unit_inst_n18), .A1(hazard_detection_unit_inst_n19), 
        .A2(hazard_detection_unit_inst_n20), .B0(
        hazard_detection_unit_inst_n21), .B1(hazard_detection_unit_inst_n22), 
        .Y(hazard_detection_unit_inst_n1) );
  INV_X0P5B_A12TS hazard_detection_unit_inst_u18 ( .A(decoding_op_src2[1]), 
        .Y(hazard_detection_unit_inst_n3) );
  INV_X0P5B_A12TS hazard_detection_unit_inst_u17 ( .A(decoding_op_src2[2]), 
        .Y(hazard_detection_unit_inst_n4) );
  INV_X0P5B_A12TS hazard_detection_unit_inst_u16 ( .A(decoding_op_src2[0]), 
        .Y(hazard_detection_unit_inst_n5) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u15 ( .A(mem_op_dest[0]), .B(
        decoding_op_src2[0]), .Y(hazard_detection_unit_inst_n11) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u14 ( .A(mem_op_dest[2]), .B(
        decoding_op_src2[2]), .Y(hazard_detection_unit_inst_n12) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u13 ( .A(mem_op_dest[1]), .B(
        decoding_op_src2[1]), .Y(hazard_detection_unit_inst_n13) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u12 ( .A(ex_op_dest[2]), .B(
        hazard_detection_unit_inst_n4), .Y(hazard_detection_unit_inst_n16) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u11 ( .A(ex_op_dest[0]), .B(
        hazard_detection_unit_inst_n5), .Y(hazard_detection_unit_inst_n17) );
  NOR2_X0P5A_A12TS hazard_detection_unit_inst_u10 ( .A(
        hazard_detection_unit_inst_n16), .B(hazard_detection_unit_inst_n17), 
        .Y(hazard_detection_unit_inst_n14) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u9 ( .A(ex_op_dest[1]), .B(
        decoding_op_src2[1]), .Y(hazard_detection_unit_inst_n15) );
  AOI32_X0P5M_A12TS hazard_detection_unit_inst_u8 ( .A0(
        hazard_detection_unit_inst_n11), .A1(hazard_detection_unit_inst_n12), 
        .A2(hazard_detection_unit_inst_n13), .B0(
        hazard_detection_unit_inst_n14), .B1(hazard_detection_unit_inst_n15), 
        .Y(hazard_detection_unit_inst_n6) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u7 ( .A(reg_write_dest[0]), .B(
        decoding_op_src2[0]), .Y(hazard_detection_unit_inst_n8) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u6 ( .A(reg_write_dest[2]), .B(
        decoding_op_src2[2]), .Y(hazard_detection_unit_inst_n9) );
  XNOR2_X0P5M_A12TS hazard_detection_unit_inst_u5 ( .A(reg_write_dest[1]), .B(
        decoding_op_src2[1]), .Y(hazard_detection_unit_inst_n10) );
  NAND3_X0P5A_A12TS hazard_detection_unit_inst_u4 ( .A(
        hazard_detection_unit_inst_n8), .B(hazard_detection_unit_inst_n9), .C(
        hazard_detection_unit_inst_n10), .Y(hazard_detection_unit_inst_n7) );
  AOI32_X0P5M_A12TS hazard_detection_unit_inst_u3 ( .A0(
        hazard_detection_unit_inst_n3), .A1(hazard_detection_unit_inst_n4), 
        .A2(hazard_detection_unit_inst_n5), .B0(hazard_detection_unit_inst_n6), 
        .B1(hazard_detection_unit_inst_n7), .Y(hazard_detection_unit_inst_n2)
         );
  NOR2_X1A_A12TS hazard_detection_unit_inst_u2 ( .A(
        hazard_detection_unit_inst_n1), .B(hazard_detection_unit_inst_n2), .Y(
        pipeline_stall_n) );
endmodule

